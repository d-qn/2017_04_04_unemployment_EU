"age","geo","time","values","geo.full"
"Y15-24","AT",2015,10.6,"Austria"
"Y15-24","AT1",2015,13.9,"Ostösterreich"
"Y15-24","AT11",2015,NA,"Burgenland (AT)"
"Y15-24","AT12",2015,10.6,"Niederösterreich"
"Y15-24","AT13",2015,18,"Wien"
"Y15-24","AT2",2015,9.8,"Südösterreich"
"Y15-24","AT21",2015,10.2,"Kärnten"
"Y15-24","AT22",2015,9.7,"Steiermark"
"Y15-24","AT3",2015,7.6,"Westösterreich"
"Y15-24","AT31",2015,9,"Oberösterreich"
"Y15-24","AT32",2015,NA,"Salzburg"
"Y15-24","AT33",2015,NA,"Tirol"
"Y15-24","AT34",2015,NA,"Vorarlberg"
"Y15-24","BE",2015,22.1,"Belgium"
"Y15-24","BE1",2015,36.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2015,36.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2015,15.2,"Vlaams Gewest"
"Y15-24","BE21",2015,15.8,"Prov. Antwerpen"
"Y15-24","BE22",2015,16.2,"Prov. Limburg (BE)"
"Y15-24","BE23",2015,16.4,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2015,17.5,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2015,10.6,"Prov. West-Vlaanderen"
"Y15-24","BE3",2015,32.2,"Région wallonne"
"Y15-24","BE31",2015,26.5,"Prov. Brabant Wallon"
"Y15-24","BE32",2015,36.7,"Prov. Hainaut"
"Y15-24","BE33",2015,30.7,"Prov. Liège"
"Y15-24","BE34",2015,19.6,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2015,35.5,"Prov. Namur"
"Y15-24","BG",2015,21.6,"Bulgaria"
"Y15-24","BG3",2015,25.8,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2015,31.7,"Severozapaden"
"Y15-24","BG32",2015,23.3,"Severen tsentralen"
"Y15-24","BG33",2015,20.5,"Severoiztochen"
"Y15-24","BG34",2015,29.7,"Yugoiztochen"
"Y15-24","BG4",2015,17.9,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2015,14.7,"Yugozapaden"
"Y15-24","BG42",2015,22.8,"Yuzhen tsentralen"
"Y15-24","CH",2015,8.6,"Switzerland"
"Y15-24","CH0",2015,8.6,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2015,16,"Région lémanique"
"Y15-24","CH02",2015,7.8,"Espace Mittelland"
"Y15-24","CH03",2015,8.6,"Nordwestschweiz"
"Y15-24","CH04",2015,5.6,"Zürich"
"Y15-24","CH05",2015,6.1,"Ostschweiz"
"Y15-24","CH06",2015,5.8,"Zentralschweiz"
"Y15-24","CH07",2015,11.5,"Ticino"
"Y15-24","CY",2015,32.8,"Cyprus"
"Y15-24","CY0",2015,32.8,"Kypros"
"Y15-24","CY00",2015,32.8,"Kypros"
"Y15-24","CZ",2015,12.6,"Czech Republic"
"Y15-24","CZ0",2015,12.6,"Ceská republika"
"Y15-24","CZ01",2015,10.6,"Praha"
"Y15-24","CZ02",2015,11.2,"Strední Cechy"
"Y15-24","CZ03",2015,8.9,"Jihozápad"
"Y15-24","CZ04",2015,17.6,"Severozápad"
"Y15-24","CZ05",2015,11.6,"Severovýchod"
"Y15-24","CZ06",2015,13.1,"Jihovýchod"
"Y15-24","CZ07",2015,10.6,"Strední Morava"
"Y15-24","CZ08",2015,16.2,"Moravskoslezsko"
"Y15-24","DE",2015,7.2,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2015,6.1,"Baden-Württemberg"
"Y15-24","DE11",2015,7,"Stuttgart"
"Y15-24","DE12",2015,5.8,"Karlsruhe"
"Y15-24","DE13",2015,4.7,"Freiburg"
"Y15-24","DE14",2015,6,"Tübingen"
"Y15-24","DE2",2015,4.2,"Bayern"
"Y15-24","DE21",2015,3.4,"Oberbayern"
"Y15-24","DE22",2015,NA,"Niederbayern"
"Y15-24","DE23",2015,NA,"Oberpfalz"
"Y15-24","DE24",2015,NA,"Oberfranken"
"Y15-24","DE25",2015,5.2,"Mittelfranken"
"Y15-24","DE26",2015,NA,"Unterfranken"
"Y15-24","DE27",2015,NA,"Schwaben"
"Y15-24","DE3",2015,15.2,"Berlin"
"Y15-24","DE30",2015,15.2,"Berlin"
"Y15-24","DE4",2015,8,"Brandenburg"
"Y15-24","DE40",2015,8,"Brandenburg"
"Y15-24","DE5",2015,NA,"Bremen"
"Y15-24","DE50",2015,NA,"Bremen"
"Y15-24","DE6",2015,7.4,"Hamburg"
"Y15-24","DE60",2015,7.4,"Hamburg"
"Y15-24","DE7",2015,6.8,"Hessen"
"Y15-24","DE71",2015,7,"Darmstadt"
"Y15-24","DE72",2015,NA,"Gießen"
"Y15-24","DE73",2015,NA,"Kassel"
"Y15-24","DE8",2015,10.7,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2015,10.7,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2015,6.4,"Niedersachsen"
"Y15-24","DE91",2015,NA,"Braunschweig"
"Y15-24","DE92",2015,7.7,"Hannover"
"Y15-24","DE93",2015,6.6,"Lüneburg"
"Y15-24","DE94",2015,5.7,"Weser-Ems"
"Y15-24","DEA",2015,8.4,"Nordrhein-Westfalen"
"Y15-24","DEA1",2015,8.9,"Düsseldorf"
"Y15-24","DEA2",2015,6.9,"Köln"
"Y15-24","DEA3",2015,8.2,"Münster"
"Y15-24","DEA4",2015,8.5,"Detmold"
"Y15-24","DEA5",2015,9.4,"Arnsberg"
"Y15-24","DEB",2015,7.4,"Rheinland-Pfalz"
"Y15-24","DEB1",2015,NA,"Koblenz"
"Y15-24","DEB2",2015,NA,"Trier"
"Y15-24","DEB3",2015,9.7,"Rheinhessen-Pfalz"
"Y15-24","DEC",2015,NA,"Saarland"
"Y15-24","DEC0",2015,NA,"Saarland"
"Y15-24","DED",2015,8.7,"Sachsen"
"Y15-24","DED2",2015,9.5,"Dresden"
"Y15-24","DED4",2015,NA,"Chemnitz"
"Y15-24","DED5",2015,NA,"Leipzig"
"Y15-24","DEE",2015,13.1,"Sachsen-Anhalt"
"Y15-24","DEE0",2015,13.1,"Sachsen-Anhalt"
"Y15-24","DEF",2015,8.2,"Schleswig-Holstein"
"Y15-24","DEF0",2015,8.2,"Schleswig-Holstein"
"Y15-24","DEG",2015,9.6,"Thüringen"
"Y15-24","DEG0",2015,9.6,"Thüringen"
"Y15-24","DK",2015,10.8,"Denmark"
"Y15-24","DK0",2015,10.8,"Danmark"
"Y15-24","DK01",2015,10,"Hovedstaden"
"Y15-24","DK02",2015,11.3,"Sjælland"
"Y15-24","DK03",2015,11.4,"Syddanmark"
"Y15-24","DK04",2015,10.4,"Midtjylland"
"Y15-24","DK05",2015,12.8,"Nordjylland"
"Y15-24","EA17",2015,22.5,"Euro area (17 countries)"
"Y15-24","EA18",2015,22.4,"Euro area (18 countries)"
"Y15-24","EA19",2015,22.4,"Euro area (19 countries)"
"Y15-24","EE",2015,13.1,"Estonia"
"Y15-24","EE0",2015,13.1,"Eesti"
"Y15-24","EE00",2015,13.1,"Eesti"
"Y15-24","EL",2015,49.8,"Greece"
"Y15-24","EL3",2015,47.2,"Attiki"
"Y15-24","EL30",2015,47.2,"Attiki"
"Y15-24","EL4",2015,38.4,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2015,42.1,"Voreio Aigaio"
"Y15-24","EL42",2015,33.8,"Notio Aigaio"
"Y15-24","EL43",2015,40.4,"Kriti"
"Y15-24","EL5",2015,52.6,"Voreia Ellada"
"Y15-24","EL51",2015,53.8,"Anatoliki Makedonia, Thraki"
"Y15-24","EL52",2015,51.9,"Kentriki Makedonia"
"Y15-24","EL53",2015,49.4,"Dytiki Makedonia"
"Y15-24","EL54",2015,58.6,"Ipeiros"
"Y15-24","EL6",2015,55.6,"Kentriki Ellada"
"Y15-24","EL61",2015,60.3,"Thessalia"
"Y15-24","EL62",2015,54.6,"Ionia Nisia"
"Y15-24","EL63",2015,54.6,"Dytiki Ellada"
"Y15-24","EL64",2015,55.4,"Sterea Ellada"
"Y15-24","EL65",2015,50.5,"Peloponnisos"
"Y15-24","ES",2015,48.3,"Spain"
"Y15-24","ES1",2015,42.7,"Noroeste (ES)"
"Y15-24","ES11",2015,43.5,"Galicia"
"Y15-24","ES12",2015,41.9,"Principado de Asturias"
"Y15-24","ES13",2015,39.6,"Cantabria"
"Y15-24","ES2",2015,40.4,"Noreste (ES)"
"Y15-24","ES21",2015,40.4,"País Vasco"
"Y15-24","ES22",2015,38.1,"Comunidad Foral de Navarra"
"Y15-24","ES23",2015,40.6,"La Rioja"
"Y15-24","ES24",2015,41.2,"Aragón"
"Y15-24","ES3",2015,44.2,"Comunidad de Madrid"
"Y15-24","ES30",2015,44.2,"Comunidad de Madrid"
"Y15-24","ES4",2015,53.5,"Centro (ES)"
"Y15-24","ES41",2015,48,"Castilla y León"
"Y15-24","ES42",2015,57.2,"Castilla-la Mancha"
"Y15-24","ES43",2015,55.4,"Extremadura"
"Y15-24","ES5",2015,44.4,"Este (ES)"
"Y15-24","ES51",2015,42.3,"Cataluña"
"Y15-24","ES52",2015,48.3,"Comunidad Valenciana"
"Y15-24","ES53",2015,42.2,"Illes Balears"
"Y15-24","ES6",2015,56.2,"Sur (ES)"
"Y15-24","ES61",2015,56.8,"Andalucía"
"Y15-24","ES62",2015,50.6,"Región de Murcia"
"Y15-24","ES63",2015,79.2,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2015,72,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2015,53.5,"Canarias (ES)"
"Y15-24","ES70",2015,53.5,"Canarias (ES)"
"Y15-24","EU15",2015,20.3,"European Union (15 countries)"
"Y15-24","EU27",2015,20.2,"European Union (27 countries)"
"Y15-24","EU28",2015,20.3,"European Union (28 countries)"
"Y15-24","FI",2015,22.4,"Finland"
"Y15-24","FI1",2015,22.5,"Manner-Suomi"
"Y15-24","FI19",2015,24.1,"Länsi-Suomi"
"Y15-24","FI1B",2015,19.1,"Helsinki-Uusimaa"
"Y15-24","FI1C",2015,22.7,"Etelä-Suomi"
"Y15-24","FI1D",2015,25.1,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2015,NA,"Åland"
"Y15-24","FI20",2015,NA,"Åland"
"Y15-24","FR",2015,24.7,"France"
"Y15-24","FR1",2015,23.2,"Île de France"
"Y15-24","FR10",2015,23.2,"Île de France"
"Y15-24","FR2",2015,23.7,"Bassin Parisien"
"Y15-24","FR21",2015,30.3,"Champagne-Ardenne"
"Y15-24","FR22",2015,22.8,"Picardie"
"Y15-24","FR23",2015,23.9,"Haute-Normandie"
"Y15-24","FR24",2015,24.5,"Centre (FR)"
"Y15-24","FR25",2015,18.7,"Basse-Normandie"
"Y15-24","FR26",2015,22.4,"Bourgogne"
"Y15-24","FR3",2015,30.1,"Nord - Pas-de-Calais"
"Y15-24","FR30",2015,30.1,"Nord - Pas-de-Calais"
"Y15-24","FR4",2015,27.1,"Est (FR)"
"Y15-24","FR41",2015,29,"Lorraine"
"Y15-24","FR42",2015,26.8,"Alsace"
"Y15-24","FR43",2015,24,"Franche-Comté"
"Y15-24","FR5",2015,22,"Ouest (FR)"
"Y15-24","FR51",2015,23.8,"Pays de la Loire"
"Y15-24","FR52",2015,18.7,"Bretagne"
"Y15-24","FR53",2015,24,"Poitou-Charentes"
"Y15-24","FR6",2015,23.5,"Sud-Ouest (FR)"
"Y15-24","FR61",2015,23.5,"Aquitaine"
"Y15-24","FR62",2015,23.4,"Midi-Pyrénées"
"Y15-24","FR63",2015,23.7,"Limousin"
"Y15-24","FR7",2015,20.3,"Centre-Est (FR)"
"Y15-24","FR71",2015,20.5,"Rhône-Alpes"
"Y15-24","FR72",2015,19.4,"Auvergne"
"Y15-24","FR8",2015,26.9,"Méditerranée"
"Y15-24","FR81",2015,31.9,"Languedoc-Roussillon"
"Y15-24","FR82",2015,24.1,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2015,NA,"Corse"
"Y15-24","FRA",2015,51.3,"Départements d'outre-mer"
"Y15-24","FRA1",2015,55.3,"Guadeloupe"
"Y15-24","FRA2",2015,47.3,"Martinique"
"Y15-24","FRA3",2015,45.4,"Guyane"
"Y15-24","FRA4",2015,51.2,"La Réunion"
"Y15-24","FRA5",2015,60.7,"Mayotte"
"Y15-24","HR",2015,42.3,"Croatia"
"Y15-24","HR0",2015,42.3,"Hrvatska"
"Y15-24","HR03",2015,43.8,"Jadranska Hrvatska"
"Y15-24","HR04",2015,41.6,"Kontinentalna Hrvatska"
"Y15-24","HU",2015,17.3,"Hungary"
"Y15-24","HU1",2015,13.2,"Közép-Magyarország"
"Y15-24","HU10",2015,13.2,"Közép-Magyarország"
"Y15-24","HU2",2015,13.2,"Dunántúl"
"Y15-24","HU21",2015,9.7,"Közép-Dunántúl"
"Y15-24","HU22",2015,12.3,"Nyugat-Dunántúl"
"Y15-24","HU23",2015,18.9,"Dél-Dunántúl"
"Y15-24","HU3",2015,22.6,"Alföld és Észak"
"Y15-24","HU31",2015,20,"Észak-Magyarország"
"Y15-24","HU32",2015,25.1,"Észak-Alföld"
"Y15-24","HU33",2015,21.9,"Dél-Alföld"
"Y15-24","IE",2015,20.9,"Ireland"
"Y15-24","IE0",2015,20.9,"Éire/Ireland"
"Y15-24","IE01",2015,24.6,"Border, Midland and Western"
"Y15-24","IE02",2015,19.6,"Southern and Eastern"
"Y15-24","IS",2015,8.8,"Iceland"
"Y15-24","IS0",2015,8.8,"Ísland"
"Y15-24","IS00",2015,8.8,"Ísland"
"Y15-24","IT",2015,40.3,"Italy"
"Y15-24","ITC",2015,34.1,"Nord-Ovest"
"Y15-24","ITC1",2015,38.1,"Piemonte"
"Y15-24","ITC2",2015,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2015,34.5,"Liguria"
"Y15-24","ITC4",2015,32.3,"Lombardia"
"Y15-24","ITF",2015,53.1,"Sud"
"Y15-24","ITF1",2015,48.1,"Abruzzo"
"Y15-24","ITF2",2015,42.7,"Molise"
"Y15-24","ITF3",2015,52.7,"Campania"
"Y15-24","ITF4",2015,51.3,"Puglia"
"Y15-24","ITF5",2015,47.7,"Basilicata"
"Y15-24","ITF6",2015,65.1,"Calabria"
"Y15-24","ITG",2015,56,"Isole"
"Y15-24","ITG1",2015,55.9,"Sicilia"
"Y15-24","ITG2",2015,56.4,"Sardegna"
"Y15-24","ITH",2015,25.9,"Nord-Est"
"Y15-24","ITH1",2015,11.9,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2015,23.6,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2015,24.6,"Veneto"
"Y15-24","ITH4",2015,28.7,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2015,29.4,"Emilia-Romagna"
"Y15-24","ITI",2015,37.7,"Centro (IT)"
"Y15-24","ITI1",2015,32.7,"Toscana"
"Y15-24","ITI2",2015,38.7,"Umbria"
"Y15-24","ITI3",2015,32,"Marche"
"Y15-24","ITI4",2015,42.6,"Lazio"
"Y15-24","LT",2015,16.3,"Lithuania"
"Y15-24","LT0",2015,16.3,"Lietuva"
"Y15-24","LT00",2015,16.3,"Lietuva"
"Y15-24","LU",2015,17.3,"Luxembourg"
"Y15-24","LU0",2015,17.3,"Luxembourg"
"Y15-24","LU00",2015,17.3,"Luxembourg"
"Y15-24","LV",2015,16.3,"Latvia"
"Y15-24","LV0",2015,16.3,"Latvija"
"Y15-24","LV00",2015,16.3,"Latvija"
"Y15-24","MK",2015,47.3,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2015,47.3,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2015,47.3,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2015,11.8,"Malta"
"Y15-24","MT0",2015,11.8,"Malta"
"Y15-24","MT00",2015,11.8,"Malta"
"Y15-24","NL",2015,11.3,"Netherlands"
"Y15-24","NL1",2015,13.9,"Noord-Nederland"
"Y15-24","NL11",2015,13.2,"Groningen"
"Y15-24","NL12",2015,15.6,"Friesland (NL)"
"Y15-24","NL13",2015,12.6,"Drenthe"
"Y15-24","NL2",2015,11,"Oost-Nederland"
"Y15-24","NL21",2015,11.5,"Overijssel"
"Y15-24","NL22",2015,10.1,"Gelderland"
"Y15-24","NL23",2015,14.5,"Flevoland"
"Y15-24","NL3",2015,11.1,"West-Nederland"
"Y15-24","NL31",2015,11,"Utrecht"
"Y15-24","NL32",2015,9.3,"Noord-Holland"
"Y15-24","NL33",2015,13,"Zuid-Holland"
"Y15-24","NL34",2015,8.1,"Zeeland"
"Y15-24","NL4",2015,10.4,"Zuid-Nederland"
"Y15-24","NL41",2015,10.5,"Noord-Brabant"
"Y15-24","NL42",2015,10.4,"Limburg (NL)"
"Y15-24","NO",2015,9.9,"Norway"
"Y15-24","NO0",2015,9.9,"Norge"
"Y15-24","NO01",2015,8.9,"Oslo og Akershus"
"Y15-24","NO02",2015,9.4,"Hedmark og Oppland"
"Y15-24","NO03",2015,11.5,"Sør-Østlandet"
"Y15-24","NO04",2015,9.4,"Agder og Rogaland"
"Y15-24","NO05",2015,9.4,"Vestlandet"
"Y15-24","NO06",2015,9.8,"Trøndelag"
"Y15-24","NO07",2015,11.3,"Nord-Norge"
"Y15-24","PL",2015,20.8,"Poland"
"Y15-24","PL1",2015,19.2,"Region Centralny"
"Y15-24","PL11",2015,20.6,"Lódzkie"
"Y15-24","PL12",2015,18.5,"Mazowieckie"
"Y15-24","PL2",2015,19.6,"Region Poludniowy"
"Y15-24","PL21",2015,20.9,"Malopolskie"
"Y15-24","PL22",2015,18.5,"Slaskie"
"Y15-24","PL3",2015,29.2,"Region Wschodni"
"Y15-24","PL31",2015,29,"Lubelskie"
"Y15-24","PL32",2015,38.4,"Podkarpackie"
"Y15-24","PL33",2015,25.8,"Swietokrzyskie"
"Y15-24","PL34",2015,18.5,"Podlaskie"
"Y15-24","PL4",2015,17.8,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2015,16.1,"Wielkopolskie"
"Y15-24","PL42",2015,23.3,"Zachodniopomorskie"
"Y15-24","PL43",2015,NA,"Lubuskie"
"Y15-24","PL5",2015,17,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2015,17.2,"Dolnoslaskie"
"Y15-24","PL52",2015,16.6,"Opolskie"
"Y15-24","PL6",2015,19.7,"Region Pólnocny"
"Y15-24","PL61",2015,18.6,"Kujawsko-Pomorskie"
"Y15-24","PL62",2015,24.1,"Warminsko-Mazurskie"
"Y15-24","PL63",2015,18.6,"Pomorskie"
"Y15-24","PT",2015,32,"Portugal"
"Y15-24","PT1",2015,31.6,"Continente"
"Y15-24","PT11",2015,32.8,"Norte"
"Y15-24","PT15",2015,29.1,"Algarve"
"Y15-24","PT16",2015,28.8,"Centro (PT)"
"Y15-24","PT17",2015,30.9,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2015,37.3,"Alentejo"
"Y15-24","PT2",2015,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2015,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2015,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2015,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2015,21.7,"Romania"
"Y15-24","RO1",2015,23.1,"Macroregiunea unu"
"Y15-24","RO11",2015,18.7,"Nord-Vest"
"Y15-24","RO12",2015,28.4,"Centru"
"Y15-24","RO2",2015,16.1,"Macroregiunea doi"
"Y15-24","RO21",2015,9.3,"Nord-Est"
"Y15-24","RO22",2015,29.3,"Sud-Est"
"Y15-24","RO3",2015,26.8,"Macroregiunea trei"
"Y15-24","RO31",2015,32.3,"Sud - Muntenia"
"Y15-24","RO32",2015,14.6,"Bucuresti - Ilfov"
"Y15-24","RO4",2015,24.1,"Macroregiunea patru"
"Y15-24","RO41",2015,27.3,"Sud-Vest Oltenia"
"Y15-24","RO42",2015,19.8,"Vest"
"Y15-24","SE",2015,20.4,"Sweden"
"Y15-24","SE1",2015,20.5,"Östra Sverige"
"Y15-24","SE11",2015,19.3,"Stockholm"
"Y15-24","SE12",2015,22.1,"Östra Mellansverige"
"Y15-24","SE2",2015,19.9,"Södra Sverige"
"Y15-24","SE21",2015,17.4,"Småland med öarna"
"Y15-24","SE22",2015,23.1,"Sydsverige"
"Y15-24","SE23",2015,18.7,"Västsverige"
"Y15-24","SE3",2015,21.4,"Norra Sverige"
"Y15-24","SE31",2015,23.3,"Norra Mellansverige"
"Y15-24","SE32",2015,20,"Mellersta Norrland"
"Y15-24","SE33",2015,19.7,"Övre Norrland"
"Y15-24","SI",2015,16.3,"Slovenia"
"Y15-24","SI0",2015,16.3,"Slovenija"
"Y15-24","SI03",2015,17,"Vzhodna Slovenija"
"Y15-24","SI04",2015,15.5,"Zahodna Slovenija"
"Y15-24","SK",2015,26.5,"Slovakia"
"Y15-24","SK0",2015,26.5,"Slovensko"
"Y15-24","SK01",2015,14.5,"Bratislavský kraj"
"Y15-24","SK02",2015,21.8,"Západné Slovensko"
"Y15-24","SK03",2015,30.5,"Stredné Slovensko"
"Y15-24","SK04",2015,31.5,"Východné Slovensko"
"Y15-24","TR",2015,18.5,"Turkey"
"Y15-24","TR1",2015,19.5,"Istanbul"
"Y15-24","TR10",2015,19.5,"Istanbul"
"Y15-24","TR2",2015,14.5,"Bati Marmara"
"Y15-24","TR21",2015,15.2,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2015,13.4,"Balikesir, Çanakkale"
"Y15-24","TR3",2015,18.1,"Ege"
"Y15-24","TR31",2015,24.8,"Izmir"
"Y15-24","TR32",2015,14.5,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2015,10.7,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2015,18.2,"Dogu Marmara"
"Y15-24","TR41",2015,15.6,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2015,20.7,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2015,18.4,"Bati Anadolu"
"Y15-24","TR51",2015,21.6,"Ankara"
"Y15-24","TR52",2015,12.9,"Konya, Karaman"
"Y15-24","TR6",2015,20.7,"Akdeniz"
"Y15-24","TR61",2015,18.9,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2015,16,"Adana, Mersin"
"Y15-24","TR63",2015,30.2,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2015,19.2,"Orta Anadolu"
"Y15-24","TR71",2015,19.6,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2015,19,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2015,14.6,"Bati Karadeniz"
"Y15-24","TR81",2015,18.9,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2015,16.2,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2015,12.7,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2015,16.3,"Dogu Karadeniz"
"Y15-24","TR90",2015,16.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2015,8,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2015,10.5,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2015,6.4,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2015,13.9,"Ortadogu Anadolu"
"Y15-24","TRB1",2015,17.5,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2015,11.8,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2015,22.6,"Güneydogu Anadolu"
"Y15-24","TRC1",2015,16.2,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2015,20.1,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2015,35.3,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2015,14.6,"United Kingdom"
"Y15-24","UKC",2015,21.2,"North East (UK)"
"Y15-24","UKC1",2015,25.1,"Tees Valley and Durham"
"Y15-24","UKC2",2015,18.4,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2015,13.4,"North West (UK)"
"Y15-24","UKD1",2015,NA,"Cumbria"
"Y15-24","UKD3",2015,15.7,"Greater Manchester"
"Y15-24","UKD4",2015,10.2,"Lancashire"
"Y15-24","UKD6",2015,10.3,"Cheshire"
"Y15-24","UKD7",2015,15.5,"Merseyside"
"Y15-24","UKE",2015,16.5,"Yorkshire and The Humber"
"Y15-24","UKE1",2015,15.3,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2015,13.2,"North Yorkshire"
"Y15-24","UKE3",2015,15.4,"South Yorkshire"
"Y15-24","UKE4",2015,18.7,"West Yorkshire"
"Y15-24","UKF",2015,11.3,"East Midlands (UK)"
"Y15-24","UKF1",2015,11,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2015,10.8,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2015,13.9,"Lincolnshire"
"Y15-24","UKG",2015,14.8,"West Midlands (UK)"
"Y15-24","UKG1",2015,10,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2015,11.3,"Shropshire and Staffordshire"
"Y15-24","UKG3",2015,19.3,"West Midlands"
"Y15-24","UKH",2015,11.9,"East of England"
"Y15-24","UKH1",2015,11.6,"East Anglia"
"Y15-24","UKH2",2015,12.4,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2015,11.8,"Essex"
"Y15-24","UKI",2015,18.7,"London"
"Y15-24","UKI3",2015,14.3,"Inner London - West"
"Y15-24","UKI4",2015,20.8,"Inner London - East"
"Y15-24","UKI5",2015,21.2,"Outer London - East and North East"
"Y15-24","UKI6",2015,14.2,"Outer London - South"
"Y15-24","UKI7",2015,18,"Outer London - West and North West"
"Y15-24","UKJ",2015,12.1,"South East (UK)"
"Y15-24","UKJ1",2015,10.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2015,11.7,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2015,11.9,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2015,14.8,"Kent"
"Y15-24","UKK",2015,11.6,"South West (UK)"
"Y15-24","UKK1",2015,10.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2015,12.1,"Dorset and Somerset"
"Y15-24","UKK3",2015,14.7,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2015,11.4,"Devon"
"Y15-24","UKL",2015,19.1,"Wales"
"Y15-24","UKL1",2015,21,"West Wales and The Valleys"
"Y15-24","UKL2",2015,16.1,"East Wales"
"Y15-24","UKM",2015,14,"Scotland"
"Y15-24","UKM2",2015,16.4,"Eastern Scotland"
"Y15-24","UKM3",2015,15.2,"South Western Scotland"
"Y15-24","UKM5",2015,8.3,"North Eastern Scotland"
"Y15-24","UKM6",2015,NA,"Highlands and Islands"
"Y15-24","UKN",2015,19.9,"Northern Ireland (UK)"
"Y15-24","UKN0",2015,19.9,"Northern Ireland (UK)"
"Y20-64","AT",2015,5.6,"Austria"
"Y20-64","AT1",2015,7.6,"Ostösterreich"
"Y20-64","AT11",2015,5.1,"Burgenland (AT)"
"Y20-64","AT12",2015,5,"Niederösterreich"
"Y20-64","AT13",2015,10.4,"Wien"
"Y20-64","AT2",2015,5,"Südösterreich"
"Y20-64","AT21",2015,6,"Kärnten"
"Y20-64","AT22",2015,4.6,"Steiermark"
"Y20-64","AT3",2015,3.5,"Westösterreich"
"Y20-64","AT31",2015,3.9,"Oberösterreich"
"Y20-64","AT32",2015,3.4,"Salzburg"
"Y20-64","AT33",2015,3,"Tirol"
"Y20-64","AT34",2015,3.4,"Vorarlberg"
"Y20-64","BE",2015,8.4,"Belgium"
"Y20-64","BE1",2015,17.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2015,17.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2015,5,"Vlaams Gewest"
"Y20-64","BE21",2015,6.1,"Prov. Antwerpen"
"Y20-64","BE22",2015,5.8,"Prov. Limburg (BE)"
"Y20-64","BE23",2015,4.2,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2015,5,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2015,4.1,"Prov. West-Vlaanderen"
"Y20-64","BE3",2015,11.7,"Région wallonne"
"Y20-64","BE31",2015,7.7,"Prov. Brabant Wallon"
"Y20-64","BE32",2015,13.1,"Prov. Hainaut"
"Y20-64","BE33",2015,12.7,"Prov. Liège"
"Y20-64","BE34",2015,9.3,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2015,10.7,"Prov. Namur"
"Y20-64","BG",2015,9.1,"Bulgaria"
"Y20-64","BG3",2015,10.6,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2015,11.9,"Severozapaden"
"Y20-64","BG32",2015,10.5,"Severen tsentralen"
"Y20-64","BG33",2015,10.2,"Severoiztochen"
"Y20-64","BG34",2015,10.2,"Yugoiztochen"
"Y20-64","BG4",2015,7.6,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2015,6.6,"Yugozapaden"
"Y20-64","BG42",2015,9.2,"Yuzhen tsentralen"
"Y20-64","CH",2015,4.4,"Switzerland"
"Y20-64","CH0",2015,4.4,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2015,6.6,"Région lémanique"
"Y20-64","CH02",2015,4.1,"Espace Mittelland"
"Y20-64","CH03",2015,3.7,"Nordwestschweiz"
"Y20-64","CH04",2015,3.9,"Zürich"
"Y20-64","CH05",2015,4,"Ostschweiz"
"Y20-64","CH06",2015,3.2,"Zentralschweiz"
"Y20-64","CH07",2015,6.4,"Ticino"
"Y20-64","CY",2015,14.9,"Cyprus"
"Y20-64","CY0",2015,14.9,"Kypros"
"Y20-64","CY00",2015,14.9,"Kypros"
"Y20-64","CZ",2015,5,"Czech Republic"
"Y20-64","CZ0",2015,5,"Ceská republika"
"Y20-64","CZ01",2015,2.8,"Praha"
"Y20-64","CZ02",2015,3.5,"Strední Cechy"
"Y20-64","CZ03",2015,3.8,"Jihozápad"
"Y20-64","CZ04",2015,7.1,"Severozápad"
"Y20-64","CZ05",2015,5.1,"Severovýchod"
"Y20-64","CZ06",2015,4.8,"Jihovýchod"
"Y20-64","CZ07",2015,5.2,"Strední Morava"
"Y20-64","CZ08",2015,8.1,"Moravskoslezsko"
"Y20-64","DE",2015,4.6,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2015,3.1,"Baden-Württemberg"
"Y20-64","DE11",2015,3.2,"Stuttgart"
"Y20-64","DE12",2015,3.3,"Karlsruhe"
"Y20-64","DE13",2015,2.5,"Freiburg"
"Y20-64","DE14",2015,2.9,"Tübingen"
"Y20-64","DE2",2015,2.9,"Bayern"
"Y20-64","DE21",2015,2.7,"Oberbayern"
"Y20-64","DE22",2015,2.6,"Niederbayern"
"Y20-64","DE23",2015,2.7,"Oberpfalz"
"Y20-64","DE24",2015,3.9,"Oberfranken"
"Y20-64","DE25",2015,3,"Mittelfranken"
"Y20-64","DE26",2015,3,"Unterfranken"
"Y20-64","DE27",2015,3,"Schwaben"
"Y20-64","DE3",2015,9.5,"Berlin"
"Y20-64","DE30",2015,9.5,"Berlin"
"Y20-64","DE4",2015,5.8,"Brandenburg"
"Y20-64","DE40",2015,5.8,"Brandenburg"
"Y20-64","DE5",2015,5.6,"Bremen"
"Y20-64","DE50",2015,5.6,"Bremen"
"Y20-64","DE6",2015,4.3,"Hamburg"
"Y20-64","DE60",2015,4.3,"Hamburg"
"Y20-64","DE7",2015,4,"Hessen"
"Y20-64","DE71",2015,4.1,"Darmstadt"
"Y20-64","DE72",2015,3.9,"Gießen"
"Y20-64","DE73",2015,3.6,"Kassel"
"Y20-64","DE8",2015,7.8,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2015,7.8,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2015,4.2,"Niedersachsen"
"Y20-64","DE91",2015,4.9,"Braunschweig"
"Y20-64","DE92",2015,4.7,"Hannover"
"Y20-64","DE93",2015,3.5,"Lüneburg"
"Y20-64","DE94",2015,3.9,"Weser-Ems"
"Y20-64","DEA",2015,5.2,"Nordrhein-Westfalen"
"Y20-64","DEA1",2015,5.9,"Düsseldorf"
"Y20-64","DEA2",2015,4.8,"Köln"
"Y20-64","DEA3",2015,4.3,"Münster"
"Y20-64","DEA4",2015,4.6,"Detmold"
"Y20-64","DEA5",2015,5.7,"Arnsberg"
"Y20-64","DEB",2015,3.6,"Rheinland-Pfalz"
"Y20-64","DEB1",2015,3.3,"Koblenz"
"Y20-64","DEB2",2015,2.9,"Trier"
"Y20-64","DEB3",2015,3.9,"Rheinhessen-Pfalz"
"Y20-64","DEC",2015,5.7,"Saarland"
"Y20-64","DEC0",2015,5.7,"Saarland"
"Y20-64","DED",2015,6.3,"Sachsen"
"Y20-64","DED2",2015,6.2,"Dresden"
"Y20-64","DED4",2015,5.5,"Chemnitz"
"Y20-64","DED5",2015,7.7,"Leipzig"
"Y20-64","DEE",2015,8,"Sachsen-Anhalt"
"Y20-64","DEE0",2015,8,"Sachsen-Anhalt"
"Y20-64","DEF",2015,4.1,"Schleswig-Holstein"
"Y20-64","DEF0",2015,4.1,"Schleswig-Holstein"
"Y20-64","DEG",2015,5.9,"Thüringen"
"Y20-64","DEG0",2015,5.9,"Thüringen"
"Y20-64","DK",2015,5.9,"Denmark"
"Y20-64","DK0",2015,5.9,"Danmark"
"Y20-64","DK01",2015,6.5,"Hovedstaden"
"Y20-64","DK02",2015,5.6,"Sjælland"
"Y20-64","DK03",2015,5.7,"Syddanmark"
"Y20-64","DK04",2015,5.4,"Midtjylland"
"Y20-64","DK05",2015,6.1,"Nordjylland"
"Y20-64","EA17",2015,10.7,"Euro area (17 countries)"
"Y20-64","EA18",2015,10.7,"Euro area (18 countries)"
"Y20-64","EA19",2015,10.7,"Euro area (19 countries)"
"Y20-64","EE",2015,6.1,"Estonia"
"Y20-64","EE0",2015,6.1,"Eesti"
"Y20-64","EE00",2015,6.1,"Eesti"
"Y20-64","EL",2015,24.9,"Greece"
"Y20-64","EL3",2015,25.1,"Attiki"
"Y20-64","EL30",2015,25.1,"Attiki"
"Y20-64","EL4",2015,20.4,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2015,17.8,"Voreio Aigaio"
"Y20-64","EL42",2015,14.6,"Notio Aigaio"
"Y20-64","EL43",2015,24.3,"Kriti"
"Y20-64","EL5",2015,25.7,"Voreia Ellada"
"Y20-64","EL51",2015,23,"Anatoliki Makedonia, Thraki"
"Y20-64","EL52",2015,26,"Kentriki Makedonia"
"Y20-64","EL53",2015,30.9,"Dytiki Makedonia"
"Y20-64","EL54",2015,24.7,"Ipeiros"
"Y20-64","EL6",2015,25.7,"Kentriki Ellada"
"Y20-64","EL61",2015,27.2,"Thessalia"
"Y20-64","EL62",2015,18.5,"Ionia Nisia"
"Y20-64","EL63",2015,28.6,"Dytiki Ellada"
"Y20-64","EL64",2015,26.1,"Sterea Ellada"
"Y20-64","EL65",2015,22.6,"Peloponnisos"
"Y20-64","ES",2015,21.7,"Spain"
"Y20-64","ES1",2015,18.9,"Noroeste (ES)"
"Y20-64","ES11",2015,19.2,"Galicia"
"Y20-64","ES12",2015,19,"Principado de Asturias"
"Y20-64","ES13",2015,17.5,"Cantabria"
"Y20-64","ES2",2015,14.9,"Noreste (ES)"
"Y20-64","ES21",2015,14.7,"País Vasco"
"Y20-64","ES22",2015,13.5,"Comunidad Foral de Navarra"
"Y20-64","ES23",2015,14.9,"La Rioja"
"Y20-64","ES24",2015,16,"Aragón"
"Y20-64","ES3",2015,16.7,"Comunidad de Madrid"
"Y20-64","ES30",2015,16.7,"Comunidad de Madrid"
"Y20-64","ES4",2015,22.9,"Centro (ES)"
"Y20-64","ES41",2015,18,"Castilla y León"
"Y20-64","ES42",2015,25.8,"Castilla-la Mancha"
"Y20-64","ES43",2015,28.6,"Extremadura"
"Y20-64","ES5",2015,19.4,"Este (ES)"
"Y20-64","ES51",2015,18.1,"Cataluña"
"Y20-64","ES52",2015,22.3,"Comunidad Valenciana"
"Y20-64","ES53",2015,16.7,"Illes Balears"
"Y20-64","ES6",2015,30.1,"Sur (ES)"
"Y20-64","ES61",2015,31.2,"Andalucía"
"Y20-64","ES62",2015,24.1,"Región de Murcia"
"Y20-64","ES63",2015,26.9,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2015,33.2,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2015,28.9,"Canarias (ES)"
"Y20-64","ES70",2015,28.9,"Canarias (ES)"
"Y20-64","EU15",2015,9.6,"European Union (15 countries)"
"Y20-64","EU27",2015,9.2,"European Union (27 countries)"
"Y20-64","EU28",2015,9.2,"European Union (28 countries)"
"Y20-64","FI",2015,8.8,"Finland"
"Y20-64","FI1",2015,8.8,"Manner-Suomi"
"Y20-64","FI19",2015,9.2,"Länsi-Suomi"
"Y20-64","FI1B",2015,7.5,"Helsinki-Uusimaa"
"Y20-64","FI1C",2015,9.5,"Etelä-Suomi"
"Y20-64","FI1D",2015,9.9,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2015,NA,"Åland"
"Y20-64","FI20",2015,NA,"Åland"
"Y20-64","FR",2015,10.1,"France"
"Y20-64","FR1",2015,9.4,"Île de France"
"Y20-64","FR10",2015,9.4,"Île de France"
"Y20-64","FR2",2015,10,"Bassin Parisien"
"Y20-64","FR21",2015,12.5,"Champagne-Ardenne"
"Y20-64","FR22",2015,10.5,"Picardie"
"Y20-64","FR23",2015,10.1,"Haute-Normandie"
"Y20-64","FR24",2015,10.4,"Centre (FR)"
"Y20-64","FR25",2015,7.9,"Basse-Normandie"
"Y20-64","FR26",2015,8.3,"Bourgogne"
"Y20-64","FR3",2015,13.7,"Nord - Pas-de-Calais"
"Y20-64","FR30",2015,13.7,"Nord - Pas-de-Calais"
"Y20-64","FR4",2015,10.1,"Est (FR)"
"Y20-64","FR41",2015,11.8,"Lorraine"
"Y20-64","FR42",2015,9,"Alsace"
"Y20-64","FR43",2015,8.6,"Franche-Comté"
"Y20-64","FR5",2015,8.3,"Ouest (FR)"
"Y20-64","FR51",2015,8.6,"Pays de la Loire"
"Y20-64","FR52",2015,7.4,"Bretagne"
"Y20-64","FR53",2015,9.3,"Poitou-Charentes"
"Y20-64","FR6",2015,8.9,"Sud-Ouest (FR)"
"Y20-64","FR61",2015,9.5,"Aquitaine"
"Y20-64","FR62",2015,8.2,"Midi-Pyrénées"
"Y20-64","FR63",2015,8.6,"Limousin"
"Y20-64","FR7",2015,8.7,"Centre-Est (FR)"
"Y20-64","FR71",2015,8.8,"Rhône-Alpes"
"Y20-64","FR72",2015,8.2,"Auvergne"
"Y20-64","FR8",2015,11.2,"Méditerranée"
"Y20-64","FR81",2015,12.5,"Languedoc-Roussillon"
"Y20-64","FR82",2015,10.7,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2015,8,"Corse"
"Y20-64","FRA",2015,22.2,"Départements d'outre-mer"
"Y20-64","FRA1",2015,23.4,"Guadeloupe"
"Y20-64","FRA2",2015,18.4,"Martinique"
"Y20-64","FRA3",2015,21.2,"Guyane"
"Y20-64","FRA4",2015,23.4,"La Réunion"
"Y20-64","FRA5",2015,23,"Mayotte"
"Y20-64","HR",2015,15.5,"Croatia"
"Y20-64","HR0",2015,15.5,"Hrvatska"
"Y20-64","HR03",2015,16.2,"Jadranska Hrvatska"
"Y20-64","HR04",2015,15.2,"Kontinentalna Hrvatska"
"Y20-64","HU",2015,6.7,"Hungary"
"Y20-64","HU1",2015,5.3,"Közép-Magyarország"
"Y20-64","HU10",2015,5.3,"Közép-Magyarország"
"Y20-64","HU2",2015,5.1,"Dunántúl"
"Y20-64","HU21",2015,4.4,"Közép-Dunántúl"
"Y20-64","HU22",2015,3.5,"Nyugat-Dunántúl"
"Y20-64","HU23",2015,7.9,"Dél-Dunántúl"
"Y20-64","HU3",2015,9,"Alföld és Észak"
"Y20-64","HU31",2015,8.4,"Észak-Magyarország"
"Y20-64","HU32",2015,10.6,"Észak-Alföld"
"Y20-64","HU33",2015,7.7,"Dél-Alföld"
"Y20-64","IE",2015,9.2,"Ireland"
"Y20-64","IE0",2015,9.2,"Éire/Ireland"
"Y20-64","IE01",2015,10.5,"Border, Midland and Western"
"Y20-64","IE02",2015,8.8,"Southern and Eastern"
"Y20-64","IS",2015,3.5,"Iceland"
"Y20-64","IS0",2015,3.5,"Ísland"
"Y20-64","IS00",2015,3.5,"Ísland"
"Y20-64","IT",2015,11.7,"Italy"
"Y20-64","ITC",2015,8.4,"Nord-Ovest"
"Y20-64","ITC1",2015,10,"Piemonte"
"Y20-64","ITC2",2015,8.7,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2015,9.2,"Liguria"
"Y20-64","ITC4",2015,7.7,"Lombardia"
"Y20-64","ITF",2015,18.6,"Sud"
"Y20-64","ITF1",2015,12.5,"Abruzzo"
"Y20-64","ITF2",2015,13.9,"Molise"
"Y20-64","ITF3",2015,19.3,"Campania"
"Y20-64","ITF4",2015,19.2,"Puglia"
"Y20-64","ITF5",2015,13.4,"Basilicata"
"Y20-64","ITF6",2015,22.7,"Calabria"
"Y20-64","ITG",2015,19.9,"Isole"
"Y20-64","ITG1",2015,21,"Sicilia"
"Y20-64","ITG2",2015,17.4,"Sardegna"
"Y20-64","ITH",2015,7.2,"Nord-Est"
"Y20-64","ITH1",2015,3.7,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2015,6.7,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2015,7.1,"Veneto"
"Y20-64","ITH4",2015,7.9,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2015,7.6,"Emilia-Romagna"
"Y20-64","ITI",2015,10.6,"Centro (IT)"
"Y20-64","ITI1",2015,9.2,"Toscana"
"Y20-64","ITI2",2015,10.3,"Umbria"
"Y20-64","ITI3",2015,9.9,"Marche"
"Y20-64","ITI4",2015,11.7,"Lazio"
"Y20-64","LT",2015,9.2,"Lithuania"
"Y20-64","LT0",2015,9.2,"Lietuva"
"Y20-64","LT00",2015,9.2,"Lietuva"
"Y20-64","LU",2015,6.3,"Luxembourg"
"Y20-64","LU0",2015,6.3,"Luxembourg"
"Y20-64","LU00",2015,6.3,"Luxembourg"
"Y20-64","LV",2015,9.9,"Latvia"
"Y20-64","LV0",2015,9.9,"Latvija"
"Y20-64","LV00",2015,9.9,"Latvija"
"Y20-64","MK",2015,26,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2015,26,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2015,26,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2015,4.9,"Malta"
"Y20-64","MT0",2015,4.9,"Malta"
"Y20-64","MT00",2015,4.9,"Malta"
"Y20-64","NL",2015,6.4,"Netherlands"
"Y20-64","NL1",2015,7.7,"Noord-Nederland"
"Y20-64","NL11",2015,8.8,"Groningen"
"Y20-64","NL12",2015,7.2,"Friesland (NL)"
"Y20-64","NL13",2015,7,"Drenthe"
"Y20-64","NL2",2015,6,"Oost-Nederland"
"Y20-64","NL21",2015,6.2,"Overijssel"
"Y20-64","NL22",2015,5.8,"Gelderland"
"Y20-64","NL23",2015,7,"Flevoland"
"Y20-64","NL3",2015,6.5,"West-Nederland"
"Y20-64","NL31",2015,6,"Utrecht"
"Y20-64","NL32",2015,5.8,"Noord-Holland"
"Y20-64","NL33",2015,7.3,"Zuid-Holland"
"Y20-64","NL34",2015,5,"Zeeland"
"Y20-64","NL4",2015,5.8,"Zuid-Nederland"
"Y20-64","NL41",2015,5.9,"Noord-Brabant"
"Y20-64","NL42",2015,5.7,"Limburg (NL)"
"Y20-64","NO",2015,4,"Norway"
"Y20-64","NO0",2015,4,"Norge"
"Y20-64","NO01",2015,4.5,"Oslo og Akershus"
"Y20-64","NO02",2015,4.2,"Hedmark og Oppland"
"Y20-64","NO03",2015,4,"Sør-Østlandet"
"Y20-64","NO04",2015,4.4,"Agder og Rogaland"
"Y20-64","NO05",2015,3.4,"Vestlandet"
"Y20-64","NO06",2015,3.5,"Trøndelag"
"Y20-64","NO07",2015,2.9,"Nord-Norge"
"Y20-64","PL",2015,7.4,"Poland"
"Y20-64","PL1",2015,6.8,"Region Centralny"
"Y20-64","PL11",2015,7.6,"Lódzkie"
"Y20-64","PL12",2015,6.4,"Mazowieckie"
"Y20-64","PL2",2015,7.1,"Region Poludniowy"
"Y20-64","PL21",2015,7.1,"Malopolskie"
"Y20-64","PL22",2015,7.1,"Slaskie"
"Y20-64","PL3",2015,9.7,"Region Wschodni"
"Y20-64","PL31",2015,9.3,"Lubelskie"
"Y20-64","PL32",2015,11.7,"Podkarpackie"
"Y20-64","PL33",2015,10,"Swietokrzyskie"
"Y20-64","PL34",2015,6.9,"Podlaskie"
"Y20-64","PL4",2015,6.2,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2015,5.7,"Wielkopolskie"
"Y20-64","PL42",2015,7.3,"Zachodniopomorskie"
"Y20-64","PL43",2015,6.4,"Lubuskie"
"Y20-64","PL5",2015,6.8,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2015,6.9,"Dolnoslaskie"
"Y20-64","PL52",2015,6.5,"Opolskie"
"Y20-64","PL6",2015,7.6,"Region Pólnocny"
"Y20-64","PL61",2015,7.8,"Kujawsko-Pomorskie"
"Y20-64","PL62",2015,9.4,"Warminsko-Mazurskie"
"Y20-64","PL63",2015,6.5,"Pomorskie"
"Y20-64","PT",2015,12.5,"Portugal"
"Y20-64","PT1",2015,12.5,"Continente"
"Y20-64","PT11",2015,13.7,"Norte"
"Y20-64","PT15",2015,12.5,"Algarve"
"Y20-64","PT16",2015,9.6,"Centro (PT)"
"Y20-64","PT17",2015,12.9,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2015,13.5,"Alentejo"
"Y20-64","PT2",2015,12.5,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2015,12.5,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2015,14.8,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2015,14.8,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2015,6.7,"Romania"
"Y20-64","RO1",2015,5.6,"Macroregiunea unu"
"Y20-64","RO11",2015,4.5,"Nord-Vest"
"Y20-64","RO12",2015,6.9,"Centru"
"Y20-64","RO2",2015,5.7,"Macroregiunea doi"
"Y20-64","RO21",2015,3.8,"Nord-Est"
"Y20-64","RO22",2015,8.6,"Sud-Est"
"Y20-64","RO3",2015,7.8,"Macroregiunea trei"
"Y20-64","RO31",2015,10.1,"Sud - Muntenia"
"Y20-64","RO32",2015,5.2,"Bucuresti - Ilfov"
"Y20-64","RO4",2015,7.9,"Macroregiunea patru"
"Y20-64","RO41",2015,10.5,"Sud-Vest Oltenia"
"Y20-64","RO42",2015,5.1,"Vest"
"Y20-64","SE",2015,6.7,"Sweden"
"Y20-64","SE1",2015,6.7,"Östra Sverige"
"Y20-64","SE11",2015,6.3,"Stockholm"
"Y20-64","SE12",2015,7.2,"Östra Mellansverige"
"Y20-64","SE2",2015,6.7,"Södra Sverige"
"Y20-64","SE21",2015,5.2,"Småland med öarna"
"Y20-64","SE22",2015,8.8,"Sydsverige"
"Y20-64","SE23",2015,5.9,"Västsverige"
"Y20-64","SE3",2015,6.7,"Norra Sverige"
"Y20-64","SE31",2015,7,"Norra Mellansverige"
"Y20-64","SE32",2015,6.6,"Mellersta Norrland"
"Y20-64","SE33",2015,6.3,"Övre Norrland"
"Y20-64","SI",2015,9,"Slovenia"
"Y20-64","SI0",2015,9,"Slovenija"
"Y20-64","SI03",2015,10.4,"Vzhodna Slovenija"
"Y20-64","SI04",2015,7.5,"Zahodna Slovenija"
"Y20-64","SK",2015,11.3,"Slovakia"
"Y20-64","SK0",2015,11.3,"Slovensko"
"Y20-64","SK01",2015,5.6,"Bratislavský kraj"
"Y20-64","SK02",2015,9.5,"Západné Slovensko"
"Y20-64","SK03",2015,12.5,"Stredné Slovensko"
"Y20-64","SK04",2015,14.7,"Východné Slovensko"
"Y20-64","TR",2015,10,"Turkey"
"Y20-64","TR1",2015,12.3,"Istanbul"
"Y20-64","TR10",2015,12.3,"Istanbul"
"Y20-64","TR2",2015,6.3,"Bati Marmara"
"Y20-64","TR21",2015,7.2,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2015,5.4,"Balikesir, Çanakkale"
"Y20-64","TR3",2015,9.2,"Ege"
"Y20-64","TR31",2015,14.5,"Izmir"
"Y20-64","TR32",2015,6.9,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2015,4,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2015,8.7,"Dogu Marmara"
"Y20-64","TR41",2015,7.7,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2015,9.7,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2015,9.5,"Bati Anadolu"
"Y20-64","TR51",2015,10.8,"Ankara"
"Y20-64","TR52",2015,6.4,"Konya, Karaman"
"Y20-64","TR6",2015,11,"Akdeniz"
"Y20-64","TR61",2015,9.2,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2015,9.8,"Adana, Mersin"
"Y20-64","TR63",2015,15.4,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2015,9.6,"Orta Anadolu"
"Y20-64","TR71",2015,9.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2015,9.4,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2015,6.9,"Bati Karadeniz"
"Y20-64","TR81",2015,7,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2015,6.9,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2015,6.8,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2015,5,"Dogu Karadeniz"
"Y20-64","TR90",2015,5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2015,4.9,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2015,5.9,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2015,4,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2015,9,"Ortadogu Anadolu"
"Y20-64","TRB1",2015,7.9,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2015,10.1,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2015,16.1,"Güneydogu Anadolu"
"Y20-64","TRC1",2015,9.4,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2015,18.1,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2015,23.2,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2015,4.6,"United Kingdom"
"Y20-64","UKC",2015,7.2,"North East (UK)"
"Y20-64","UKC1",2015,7.4,"Tees Valley and Durham"
"Y20-64","UKC2",2015,7.1,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2015,4.7,"North West (UK)"
"Y20-64","UKD1",2015,3.9,"Cumbria"
"Y20-64","UKD3",2015,5.4,"Greater Manchester"
"Y20-64","UKD4",2015,4.1,"Lancashire"
"Y20-64","UKD6",2015,3.2,"Cheshire"
"Y20-64","UKD7",2015,5.2,"Merseyside"
"Y20-64","UKE",2015,5.4,"Yorkshire and The Humber"
"Y20-64","UKE1",2015,5.8,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2015,2.4,"North Yorkshire"
"Y20-64","UKE3",2015,6.7,"South Yorkshire"
"Y20-64","UKE4",2015,5.6,"West Yorkshire"
"Y20-64","UKF",2015,4,"East Midlands (UK)"
"Y20-64","UKF1",2015,4.3,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2015,3.8,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2015,3.5,"Lincolnshire"
"Y20-64","UKG",2015,5.3,"West Midlands (UK)"
"Y20-64","UKG1",2015,2.9,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2015,4,"Shropshire and Staffordshire"
"Y20-64","UKG3",2015,7.4,"West Midlands"
"Y20-64","UKH",2015,3.5,"East of England"
"Y20-64","UKH1",2015,3.6,"East Anglia"
"Y20-64","UKH2",2015,3.4,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2015,3.6,"Essex"
"Y20-64","UKI",2015,5.5,"London"
"Y20-64","UKI3",2015,5.3,"Inner London - West"
"Y20-64","UKI4",2015,6.4,"Inner London - East"
"Y20-64","UKI5",2015,6.4,"Outer London - East and North East"
"Y20-64","UKI6",2015,4,"Outer London - South"
"Y20-64","UKI7",2015,4.7,"Outer London - West and North West"
"Y20-64","UKJ",2015,3.5,"South East (UK)"
"Y20-64","UKJ1",2015,3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2015,3.2,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2015,3.6,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2015,4.8,"Kent"
"Y20-64","UKK",2015,3.2,"South West (UK)"
"Y20-64","UKK1",2015,3.2,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2015,3.1,"Dorset and Somerset"
"Y20-64","UKK3",2015,3.5,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2015,3.2,"Devon"
"Y20-64","UKL",2015,5,"Wales"
"Y20-64","UKL1",2015,5.7,"West Wales and The Valleys"
"Y20-64","UKL2",2015,3.7,"East Wales"
"Y20-64","UKM",2015,4.9,"Scotland"
"Y20-64","UKM2",2015,5,"Eastern Scotland"
"Y20-64","UKM3",2015,5.9,"South Western Scotland"
"Y20-64","UKM5",2015,2.1,"North Eastern Scotland"
"Y20-64","UKM6",2015,3.7,"Highlands and Islands"
"Y20-64","UKN",2015,5.8,"Northern Ireland (UK)"
"Y20-64","UKN0",2015,5.8,"Northern Ireland (UK)"
"Y_GE15","AT",2015,5.7,"Austria"
"Y_GE15","AT1",2015,7.8,"Ostösterreich"
"Y_GE15","AT11",2015,5.2,"Burgenland (AT)"
"Y_GE15","AT12",2015,5.2,"Niederösterreich"
"Y_GE15","AT13",2015,10.6,"Wien"
"Y_GE15","AT2",2015,5.1,"Südösterreich"
"Y_GE15","AT21",2015,6.1,"Kärnten"
"Y_GE15","AT22",2015,4.7,"Steiermark"
"Y_GE15","AT3",2015,3.7,"Westösterreich"
"Y_GE15","AT31",2015,4.1,"Oberösterreich"
"Y_GE15","AT32",2015,3.5,"Salzburg"
"Y_GE15","AT33",2015,3,"Tirol"
"Y_GE15","AT34",2015,3.5,"Vorarlberg"
"Y_GE15","BE",2015,8.5,"Belgium"
"Y_GE15","BE1",2015,17.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2015,17.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2015,5.2,"Vlaams Gewest"
"Y_GE15","BE21",2015,6.1,"Prov. Antwerpen"
"Y_GE15","BE22",2015,6,"Prov. Limburg (BE)"
"Y_GE15","BE23",2015,4.4,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2015,5.1,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2015,4.2,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2015,11.9,"Région wallonne"
"Y_GE15","BE31",2015,7.8,"Prov. Brabant Wallon"
"Y_GE15","BE32",2015,13.3,"Prov. Hainaut"
"Y_GE15","BE33",2015,12.8,"Prov. Liège"
"Y_GE15","BE34",2015,9.3,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2015,10.9,"Prov. Namur"
"Y_GE15","BG",2015,9.1,"Bulgaria"
"Y_GE15","BG3",2015,10.7,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2015,12.1,"Severozapaden"
"Y_GE15","BG32",2015,10.6,"Severen tsentralen"
"Y_GE15","BG33",2015,10.3,"Severoiztochen"
"Y_GE15","BG34",2015,10.4,"Yugoiztochen"
"Y_GE15","BG4",2015,7.7,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2015,6.7,"Yugozapaden"
"Y_GE15","BG42",2015,9.2,"Yuzhen tsentralen"
"Y_GE15","CH",2015,4.5,"Switzerland"
"Y_GE15","CH0",2015,4.5,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2015,7,"Région lémanique"
"Y_GE15","CH02",2015,4.1,"Espace Mittelland"
"Y_GE15","CH03",2015,4,"Nordwestschweiz"
"Y_GE15","CH04",2015,3.9,"Zürich"
"Y_GE15","CH05",2015,3.8,"Ostschweiz"
"Y_GE15","CH06",2015,3.3,"Zentralschweiz"
"Y_GE15","CH07",2015,6.4,"Ticino"
"Y_GE15","CY",2015,14.9,"Cyprus"
"Y_GE15","CY0",2015,14.9,"Kypros"
"Y_GE15","CY00",2015,14.9,"Kypros"
"Y_GE15","CZ",2015,5,"Czech Republic"
"Y_GE15","CZ0",2015,5,"Ceská republika"
"Y_GE15","CZ01",2015,2.8,"Praha"
"Y_GE15","CZ02",2015,3.5,"Strední Cechy"
"Y_GE15","CZ03",2015,3.9,"Jihozápad"
"Y_GE15","CZ04",2015,7.3,"Severozápad"
"Y_GE15","CZ05",2015,5.2,"Severovýchod"
"Y_GE15","CZ06",2015,4.9,"Jihovýchod"
"Y_GE15","CZ07",2015,5.3,"Strední Morava"
"Y_GE15","CZ08",2015,8.1,"Moravskoslezsko"
"Y_GE15","DE",2015,4.6,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2015,3.1,"Baden-Württemberg"
"Y_GE15","DE11",2015,3.3,"Stuttgart"
"Y_GE15","DE12",2015,3.3,"Karlsruhe"
"Y_GE15","DE13",2015,2.5,"Freiburg"
"Y_GE15","DE14",2015,3,"Tübingen"
"Y_GE15","DE2",2015,2.9,"Bayern"
"Y_GE15","DE21",2015,2.7,"Oberbayern"
"Y_GE15","DE22",2015,2.5,"Niederbayern"
"Y_GE15","DE23",2015,2.7,"Oberpfalz"
"Y_GE15","DE24",2015,3.8,"Oberfranken"
"Y_GE15","DE25",2015,3,"Mittelfranken"
"Y_GE15","DE26",2015,3,"Unterfranken"
"Y_GE15","DE27",2015,3,"Schwaben"
"Y_GE15","DE3",2015,9.4,"Berlin"
"Y_GE15","DE30",2015,9.4,"Berlin"
"Y_GE15","DE4",2015,5.7,"Brandenburg"
"Y_GE15","DE40",2015,5.7,"Brandenburg"
"Y_GE15","DE5",2015,5.6,"Bremen"
"Y_GE15","DE50",2015,5.6,"Bremen"
"Y_GE15","DE6",2015,4.3,"Hamburg"
"Y_GE15","DE60",2015,4.3,"Hamburg"
"Y_GE15","DE7",2015,4,"Hessen"
"Y_GE15","DE71",2015,4.1,"Darmstadt"
"Y_GE15","DE72",2015,3.8,"Gießen"
"Y_GE15","DE73",2015,3.6,"Kassel"
"Y_GE15","DE8",2015,7.8,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2015,7.8,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2015,4.3,"Niedersachsen"
"Y_GE15","DE91",2015,4.9,"Braunschweig"
"Y_GE15","DE92",2015,4.7,"Hannover"
"Y_GE15","DE93",2015,3.5,"Lüneburg"
"Y_GE15","DE94",2015,3.9,"Weser-Ems"
"Y_GE15","DEA",2015,5.2,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2015,5.9,"Düsseldorf"
"Y_GE15","DEA2",2015,4.8,"Köln"
"Y_GE15","DEA3",2015,4.4,"Münster"
"Y_GE15","DEA4",2015,4.7,"Detmold"
"Y_GE15","DEA5",2015,5.7,"Arnsberg"
"Y_GE15","DEB",2015,3.7,"Rheinland-Pfalz"
"Y_GE15","DEB1",2015,3.4,"Koblenz"
"Y_GE15","DEB2",2015,2.9,"Trier"
"Y_GE15","DEB3",2015,4.1,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2015,5.6,"Saarland"
"Y_GE15","DEC0",2015,5.6,"Saarland"
"Y_GE15","DED",2015,6.3,"Sachsen"
"Y_GE15","DED2",2015,6.2,"Dresden"
"Y_GE15","DED4",2015,5.4,"Chemnitz"
"Y_GE15","DED5",2015,7.7,"Leipzig"
"Y_GE15","DEE",2015,8,"Sachsen-Anhalt"
"Y_GE15","DEE0",2015,8,"Sachsen-Anhalt"
"Y_GE15","DEF",2015,4.2,"Schleswig-Holstein"
"Y_GE15","DEF0",2015,4.2,"Schleswig-Holstein"
"Y_GE15","DEG",2015,5.8,"Thüringen"
"Y_GE15","DEG0",2015,5.8,"Thüringen"
"Y_GE15","DK",2015,6.2,"Denmark"
"Y_GE15","DK0",2015,6.2,"Danmark"
"Y_GE15","DK01",2015,6.7,"Hovedstaden"
"Y_GE15","DK02",2015,5.9,"Sjælland"
"Y_GE15","DK03",2015,6.1,"Syddanmark"
"Y_GE15","DK04",2015,5.6,"Midtjylland"
"Y_GE15","DK05",2015,6.3,"Nordjylland"
"Y_GE15","EA17",2015,10.9,"Euro area (17 countries)"
"Y_GE15","EA18",2015,10.9,"Euro area (18 countries)"
"Y_GE15","EA19",2015,10.8,"Euro area (19 countries)"
"Y_GE15","EE",2015,6.2,"Estonia"
"Y_GE15","EE0",2015,6.2,"Eesti"
"Y_GE15","EE00",2015,6.2,"Eesti"
"Y_GE15","EL",2015,24.9,"Greece"
"Y_GE15","EL3",2015,25.2,"Attiki"
"Y_GE15","EL30",2015,25.2,"Attiki"
"Y_GE15","EL4",2015,20.4,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2015,18,"Voreio Aigaio"
"Y_GE15","EL42",2015,14.9,"Notio Aigaio"
"Y_GE15","EL43",2015,24.2,"Kriti"
"Y_GE15","EL5",2015,25.7,"Voreia Ellada"
"Y_GE15","EL51",2015,23.4,"Anatoliki Makedonia, Thraki"
"Y_GE15","EL52",2015,26,"Kentriki Makedonia"
"Y_GE15","EL53",2015,30.7,"Dytiki Makedonia"
"Y_GE15","EL54",2015,24.5,"Ipeiros"
"Y_GE15","EL6",2015,25.5,"Kentriki Ellada"
"Y_GE15","EL61",2015,26.9,"Thessalia"
"Y_GE15","EL62",2015,19,"Ionia Nisia"
"Y_GE15","EL63",2015,28.5,"Dytiki Ellada"
"Y_GE15","EL64",2015,25.8,"Sterea Ellada"
"Y_GE15","EL65",2015,22.3,"Peloponnisos"
"Y_GE15","ES",2015,22.1,"Spain"
"Y_GE15","ES1",2015,19,"Noroeste (ES)"
"Y_GE15","ES11",2015,19.3,"Galicia"
"Y_GE15","ES12",2015,19.1,"Principado de Asturias"
"Y_GE15","ES13",2015,17.6,"Cantabria"
"Y_GE15","ES2",2015,15.1,"Noreste (ES)"
"Y_GE15","ES21",2015,14.8,"País Vasco"
"Y_GE15","ES22",2015,13.8,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2015,15.4,"La Rioja"
"Y_GE15","ES24",2015,16.3,"Aragón"
"Y_GE15","ES3",2015,17.1,"Comunidad de Madrid"
"Y_GE15","ES30",2015,17.1,"Comunidad de Madrid"
"Y_GE15","ES4",2015,23.4,"Centro (ES)"
"Y_GE15","ES41",2015,18.3,"Castilla y León"
"Y_GE15","ES42",2015,26.3,"Castilla-la Mancha"
"Y_GE15","ES43",2015,29.1,"Extremadura"
"Y_GE15","ES5",2015,20,"Este (ES)"
"Y_GE15","ES51",2015,18.6,"Cataluña"
"Y_GE15","ES52",2015,22.8,"Comunidad Valenciana"
"Y_GE15","ES53",2015,17.3,"Illes Balears"
"Y_GE15","ES6",2015,30.5,"Sur (ES)"
"Y_GE15","ES61",2015,31.5,"Andalucía"
"Y_GE15","ES62",2015,24.6,"Región de Murcia"
"Y_GE15","ES63",2015,27.6,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2015,34,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2015,29.1,"Canarias (ES)"
"Y_GE15","ES70",2015,29.1,"Canarias (ES)"
"Y_GE15","EU15",2015,9.8,"European Union (15 countries)"
"Y_GE15","EU27",2015,9.3,"European Union (27 countries)"
"Y_GE15","EU28",2015,9.4,"European Union (28 countries)"
"Y_GE15","FI",2015,9.4,"Finland"
"Y_GE15","FI1",2015,9.4,"Manner-Suomi"
"Y_GE15","FI19",2015,9.8,"Länsi-Suomi"
"Y_GE15","FI1B",2015,8,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2015,10,"Etelä-Suomi"
"Y_GE15","FI1D",2015,10.4,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2015,NA,"Åland"
"Y_GE15","FI20",2015,NA,"Åland"
"Y_GE15","FR",2015,10.4,"France"
"Y_GE15","FR1",2015,9.6,"Île de France"
"Y_GE15","FR10",2015,9.6,"Île de France"
"Y_GE15","FR2",2015,10.3,"Bassin Parisien"
"Y_GE15","FR21",2015,13,"Champagne-Ardenne"
"Y_GE15","FR22",2015,10.8,"Picardie"
"Y_GE15","FR23",2015,10.6,"Haute-Normandie"
"Y_GE15","FR24",2015,10.7,"Centre (FR)"
"Y_GE15","FR25",2015,8.2,"Basse-Normandie"
"Y_GE15","FR26",2015,8.7,"Bourgogne"
"Y_GE15","FR3",2015,14,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2015,14,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2015,10.5,"Est (FR)"
"Y_GE15","FR41",2015,12.2,"Lorraine"
"Y_GE15","FR42",2015,9.3,"Alsace"
"Y_GE15","FR43",2015,9.2,"Franche-Comté"
"Y_GE15","FR5",2015,8.7,"Ouest (FR)"
"Y_GE15","FR51",2015,9.1,"Pays de la Loire"
"Y_GE15","FR52",2015,7.8,"Bretagne"
"Y_GE15","FR53",2015,9.7,"Poitou-Charentes"
"Y_GE15","FR6",2015,9.2,"Sud-Ouest (FR)"
"Y_GE15","FR61",2015,9.8,"Aquitaine"
"Y_GE15","FR62",2015,8.5,"Midi-Pyrénées"
"Y_GE15","FR63",2015,8.9,"Limousin"
"Y_GE15","FR7",2015,9,"Centre-Est (FR)"
"Y_GE15","FR71",2015,9.1,"Rhône-Alpes"
"Y_GE15","FR72",2015,8.6,"Auvergne"
"Y_GE15","FR8",2015,11.6,"Méditerranée"
"Y_GE15","FR81",2015,12.9,"Languedoc-Roussillon"
"Y_GE15","FR82",2015,11,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2015,8.5,"Corse"
"Y_GE15","FRA",2015,22.7,"Départements d'outre-mer"
"Y_GE15","FRA1",2015,23.7,"Guadeloupe"
"Y_GE15","FRA2",2015,18.6,"Martinique"
"Y_GE15","FRA3",2015,21.9,"Guyane"
"Y_GE15","FRA4",2015,24.1,"La Réunion"
"Y_GE15","FRA5",2015,23.7,"Mayotte"
"Y_GE15","HR",2015,16.2,"Croatia"
"Y_GE15","HR0",2015,16.2,"Hrvatska"
"Y_GE15","HR03",2015,16.8,"Jadranska Hrvatska"
"Y_GE15","HR04",2015,15.9,"Kontinentalna Hrvatska"
"Y_GE15","HU",2015,6.8,"Hungary"
"Y_GE15","HU1",2015,5.3,"Közép-Magyarország"
"Y_GE15","HU10",2015,5.3,"Közép-Magyarország"
"Y_GE15","HU2",2015,5.3,"Dunántúl"
"Y_GE15","HU21",2015,4.4,"Közép-Dunántúl"
"Y_GE15","HU22",2015,3.8,"Nyugat-Dunántúl"
"Y_GE15","HU23",2015,8.1,"Dél-Dunántúl"
"Y_GE15","HU3",2015,9.2,"Alföld és Észak"
"Y_GE15","HU31",2015,8.7,"Észak-Magyarország"
"Y_GE15","HU32",2015,10.9,"Észak-Alföld"
"Y_GE15","HU33",2015,7.9,"Dél-Alföld"
"Y_GE15","IE",2015,9.4,"Ireland"
"Y_GE15","IE0",2015,9.4,"Éire/Ireland"
"Y_GE15","IE01",2015,10.6,"Border, Midland and Western"
"Y_GE15","IE02",2015,9,"Southern and Eastern"
"Y_GE15","IS",2015,4,"Iceland"
"Y_GE15","IS0",2015,4,"Ísland"
"Y_GE15","IS00",2015,4,"Ísland"
"Y_GE15","IT",2015,11.9,"Italy"
"Y_GE15","ITC",2015,8.6,"Nord-Ovest"
"Y_GE15","ITC1",2015,10.2,"Piemonte"
"Y_GE15","ITC2",2015,8.9,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2015,9.2,"Liguria"
"Y_GE15","ITC4",2015,7.9,"Lombardia"
"Y_GE15","ITF",2015,19,"Sud"
"Y_GE15","ITF1",2015,12.6,"Abruzzo"
"Y_GE15","ITF2",2015,14.3,"Molise"
"Y_GE15","ITF3",2015,19.8,"Campania"
"Y_GE15","ITF4",2015,19.7,"Puglia"
"Y_GE15","ITF5",2015,13.7,"Basilicata"
"Y_GE15","ITF6",2015,22.9,"Calabria"
"Y_GE15","ITG",2015,20.3,"Isole"
"Y_GE15","ITG1",2015,21.4,"Sicilia"
"Y_GE15","ITG2",2015,17.4,"Sardegna"
"Y_GE15","ITH",2015,7.3,"Nord-Est"
"Y_GE15","ITH1",2015,3.8,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2015,6.8,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2015,7.1,"Veneto"
"Y_GE15","ITH4",2015,8,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2015,7.7,"Emilia-Romagna"
"Y_GE15","ITI",2015,10.6,"Centro (IT)"
"Y_GE15","ITI1",2015,9.2,"Toscana"
"Y_GE15","ITI2",2015,10.4,"Umbria"
"Y_GE15","ITI3",2015,9.9,"Marche"
"Y_GE15","ITI4",2015,11.8,"Lazio"
"Y_GE15","LT",2015,9.1,"Lithuania"
"Y_GE15","LT0",2015,9.1,"Lietuva"
"Y_GE15","LT00",2015,9.1,"Lietuva"
"Y_GE15","LU",2015,6.7,"Luxembourg"
"Y_GE15","LU0",2015,6.7,"Luxembourg"
"Y_GE15","LU00",2015,6.7,"Luxembourg"
"Y_GE15","LV",2015,9.9,"Latvia"
"Y_GE15","LV0",2015,9.9,"Latvija"
"Y_GE15","LV00",2015,9.9,"Latvija"
"Y_GE15","MK",2015,26.1,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2015,26.1,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2015,26.1,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2015,5.4,"Malta"
"Y_GE15","MT0",2015,5.4,"Malta"
"Y_GE15","MT00",2015,5.4,"Malta"
"Y_GE15","NL",2015,6.9,"Netherlands"
"Y_GE15","NL1",2015,8.2,"Noord-Nederland"
"Y_GE15","NL11",2015,9.1,"Groningen"
"Y_GE15","NL12",2015,7.9,"Friesland (NL)"
"Y_GE15","NL13",2015,7.5,"Drenthe"
"Y_GE15","NL2",2015,6.6,"Oost-Nederland"
"Y_GE15","NL21",2015,6.9,"Overijssel"
"Y_GE15","NL22",2015,6.3,"Gelderland"
"Y_GE15","NL23",2015,7.9,"Flevoland"
"Y_GE15","NL3",2015,6.9,"West-Nederland"
"Y_GE15","NL31",2015,6.4,"Utrecht"
"Y_GE15","NL32",2015,6.2,"Noord-Holland"
"Y_GE15","NL33",2015,7.8,"Zuid-Holland"
"Y_GE15","NL34",2015,5.3,"Zeeland"
"Y_GE15","NL4",2015,6.4,"Zuid-Nederland"
"Y_GE15","NL41",2015,6.5,"Noord-Brabant"
"Y_GE15","NL42",2015,6.3,"Limburg (NL)"
"Y_GE15","NO",2015,4.3,"Norway"
"Y_GE15","NO0",2015,4.3,"Norge"
"Y_GE15","NO01",2015,4.7,"Oslo og Akershus"
"Y_GE15","NO02",2015,4.5,"Hedmark og Oppland"
"Y_GE15","NO03",2015,4.5,"Sør-Østlandet"
"Y_GE15","NO04",2015,4.6,"Agder og Rogaland"
"Y_GE15","NO05",2015,3.9,"Vestlandet"
"Y_GE15","NO06",2015,3.7,"Trøndelag"
"Y_GE15","NO07",2015,3.4,"Nord-Norge"
"Y_GE15","PL",2015,7.5,"Poland"
"Y_GE15","PL1",2015,6.8,"Region Centralny"
"Y_GE15","PL11",2015,7.7,"Lódzkie"
"Y_GE15","PL12",2015,6.4,"Mazowieckie"
"Y_GE15","PL2",2015,7.2,"Region Poludniowy"
"Y_GE15","PL21",2015,7.1,"Malopolskie"
"Y_GE15","PL22",2015,7.2,"Slaskie"
"Y_GE15","PL3",2015,9.7,"Region Wschodni"
"Y_GE15","PL31",2015,9.3,"Lubelskie"
"Y_GE15","PL32",2015,11.6,"Podkarpackie"
"Y_GE15","PL33",2015,10.1,"Swietokrzyskie"
"Y_GE15","PL34",2015,7,"Podlaskie"
"Y_GE15","PL4",2015,6.3,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2015,5.8,"Wielkopolskie"
"Y_GE15","PL42",2015,7.5,"Zachodniopomorskie"
"Y_GE15","PL43",2015,6.4,"Lubuskie"
"Y_GE15","PL5",2015,6.9,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2015,7,"Dolnoslaskie"
"Y_GE15","PL52",2015,6.5,"Opolskie"
"Y_GE15","PL6",2015,7.7,"Region Pólnocny"
"Y_GE15","PL61",2015,7.9,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2015,9.5,"Warminsko-Mazurskie"
"Y_GE15","PL63",2015,6.6,"Pomorskie"
"Y_GE15","PT",2015,12.4,"Portugal"
"Y_GE15","PT1",2015,12.4,"Continente"
"Y_GE15","PT11",2015,13.7,"Norte"
"Y_GE15","PT15",2015,12.5,"Algarve"
"Y_GE15","PT16",2015,9.2,"Centro (PT)"
"Y_GE15","PT17",2015,13.1,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2015,13.3,"Alentejo"
"Y_GE15","PT2",2015,12.8,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2015,12.8,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2015,14.7,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2015,14.7,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2015,6.8,"Romania"
"Y_GE15","RO1",2015,5.9,"Macroregiunea unu"
"Y_GE15","RO11",2015,4.6,"Nord-Vest"
"Y_GE15","RO12",2015,7.4,"Centru"
"Y_GE15","RO2",2015,5.8,"Macroregiunea doi"
"Y_GE15","RO21",2015,3.6,"Nord-Est"
"Y_GE15","RO22",2015,9,"Sud-Est"
"Y_GE15","RO3",2015,8,"Macroregiunea trei"
"Y_GE15","RO31",2015,10.3,"Sud - Muntenia"
"Y_GE15","RO32",2015,5.3,"Bucuresti - Ilfov"
"Y_GE15","RO4",2015,7.9,"Macroregiunea patru"
"Y_GE15","RO41",2015,10.1,"Sud-Vest Oltenia"
"Y_GE15","RO42",2015,5.4,"Vest"
"Y_GE15","SE",2015,7.4,"Sweden"
"Y_GE15","SE1",2015,7.4,"Östra Sverige"
"Y_GE15","SE11",2015,7,"Stockholm"
"Y_GE15","SE12",2015,7.9,"Östra Mellansverige"
"Y_GE15","SE2",2015,7.4,"Södra Sverige"
"Y_GE15","SE21",2015,6,"Småland med öarna"
"Y_GE15","SE22",2015,9.5,"Sydsverige"
"Y_GE15","SE23",2015,6.6,"Västsverige"
"Y_GE15","SE3",2015,7.5,"Norra Sverige"
"Y_GE15","SE31",2015,7.9,"Norra Mellansverige"
"Y_GE15","SE32",2015,7.1,"Mellersta Norrland"
"Y_GE15","SE33",2015,7.2,"Övre Norrland"
"Y_GE15","SI",2015,9,"Slovenia"
"Y_GE15","SI0",2015,9,"Slovenija"
"Y_GE15","SI03",2015,10.3,"Vzhodna Slovenija"
"Y_GE15","SI04",2015,7.5,"Zahodna Slovenija"
"Y_GE15","SK",2015,11.5,"Slovakia"
"Y_GE15","SK0",2015,11.5,"Slovensko"
"Y_GE15","SK01",2015,5.7,"Bratislavský kraj"
"Y_GE15","SK02",2015,9.7,"Západné Slovensko"
"Y_GE15","SK03",2015,12.8,"Stredné Slovensko"
"Y_GE15","SK04",2015,15,"Východné Slovensko"
"Y_GE15","TR",2015,10.2,"Turkey"
"Y_GE15","TR1",2015,12.8,"Istanbul"
"Y_GE15","TR10",2015,12.8,"Istanbul"
"Y_GE15","TR2",2015,6.4,"Bati Marmara"
"Y_GE15","TR21",2015,7.3,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2015,5.3,"Balikesir, Çanakkale"
"Y_GE15","TR3",2015,9.4,"Ege"
"Y_GE15","TR31",2015,14.9,"Izmir"
"Y_GE15","TR32",2015,6.8,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2015,4.1,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2015,8.9,"Dogu Marmara"
"Y_GE15","TR41",2015,7.7,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2015,10.1,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2015,9.7,"Bati Anadolu"
"Y_GE15","TR51",2015,11.1,"Ankara"
"Y_GE15","TR52",2015,6.5,"Konya, Karaman"
"Y_GE15","TR6",2015,11.3,"Akdeniz"
"Y_GE15","TR61",2015,9.4,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2015,9.8,"Adana, Mersin"
"Y_GE15","TR63",2015,16.3,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2015,9.8,"Orta Anadolu"
"Y_GE15","TR71",2015,9.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2015,9.7,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2015,6.7,"Bati Karadeniz"
"Y_GE15","TR81",2015,6.9,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2015,6.8,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2015,6.6,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2015,4.8,"Dogu Karadeniz"
"Y_GE15","TR90",2015,4.8,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2015,4.9,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2015,6,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2015,3.9,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2015,8.8,"Ortadogu Anadolu"
"Y_GE15","TRB1",2015,7.9,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2015,9.7,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2015,16.3,"Güneydogu Anadolu"
"Y_GE15","TRC1",2015,9.7,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2015,17.4,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2015,24.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2015,5.3,"United Kingdom"
"Y_GE15","UKC",2015,8,"North East (UK)"
"Y_GE15","UKC1",2015,8.5,"Tees Valley and Durham"
"Y_GE15","UKC2",2015,7.7,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2015,5.4,"North West (UK)"
"Y_GE15","UKD1",2015,4.2,"Cumbria"
"Y_GE15","UKD3",2015,6.5,"Greater Manchester"
"Y_GE15","UKD4",2015,4.5,"Lancashire"
"Y_GE15","UKD6",2015,3.5,"Cheshire"
"Y_GE15","UKD7",2015,5.8,"Merseyside"
"Y_GE15","UKE",2015,6.2,"Yorkshire and The Humber"
"Y_GE15","UKE1",2015,6.4,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2015,3.2,"North Yorkshire"
"Y_GE15","UKE3",2015,7.4,"South Yorkshire"
"Y_GE15","UKE4",2015,6.6,"West Yorkshire"
"Y_GE15","UKF",2015,4.6,"East Midlands (UK)"
"Y_GE15","UKF1",2015,4.8,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2015,4.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2015,4.5,"Lincolnshire"
"Y_GE15","UKG",2015,5.8,"West Midlands (UK)"
"Y_GE15","UKG1",2015,3.2,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2015,4.6,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2015,7.9,"West Midlands"
"Y_GE15","UKH",2015,4.2,"East of England"
"Y_GE15","UKH1",2015,4.3,"East Anglia"
"Y_GE15","UKH2",2015,3.8,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2015,4.3,"Essex"
"Y_GE15","UKI",2015,6.2,"London"
"Y_GE15","UKI3",2015,5.4,"Inner London - West"
"Y_GE15","UKI4",2015,7.2,"Inner London - East"
"Y_GE15","UKI5",2015,7.5,"Outer London - East and North East"
"Y_GE15","UKI6",2015,4.6,"Outer London - South"
"Y_GE15","UKI7",2015,5.5,"Outer London - West and North West"
"Y_GE15","UKJ",2015,4,"South East (UK)"
"Y_GE15","UKJ1",2015,3.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2015,3.7,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2015,4.1,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2015,5.3,"Kent"
"Y_GE15","UKK",2015,3.9,"South West (UK)"
"Y_GE15","UKK1",2015,3.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2015,3.9,"Dorset and Somerset"
"Y_GE15","UKK3",2015,4.5,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2015,3.7,"Devon"
"Y_GE15","UKL",2015,5.9,"Wales"
"Y_GE15","UKL1",2015,6.5,"West Wales and The Valleys"
"Y_GE15","UKL2",2015,4.8,"East Wales"
"Y_GE15","UKM",2015,5.7,"Scotland"
"Y_GE15","UKM2",2015,6,"Eastern Scotland"
"Y_GE15","UKM3",2015,6.6,"South Western Scotland"
"Y_GE15","UKM5",2015,3.2,"North Eastern Scotland"
"Y_GE15","UKM6",2015,4.1,"Highlands and Islands"
"Y_GE15","UKN",2015,6.1,"Northern Ireland (UK)"
"Y_GE15","UKN0",2015,6.1,"Northern Ireland (UK)"
"Y_GE25","AT",2015,5,"Austria"
"Y_GE25","AT1",2015,6.9,"Ostösterreich"
"Y_GE25","AT11",2015,4.9,"Burgenland (AT)"
"Y_GE25","AT12",2015,4.4,"Niederösterreich"
"Y_GE25","AT13",2015,9.6,"Wien"
"Y_GE25","AT2",2015,4.5,"Südösterreich"
"Y_GE25","AT21",2015,5.5,"Kärnten"
"Y_GE25","AT22",2015,4,"Steiermark"
"Y_GE25","AT3",2015,3.1,"Westösterreich"
"Y_GE25","AT31",2015,3.3,"Oberösterreich"
"Y_GE25","AT32",2015,3,"Salzburg"
"Y_GE25","AT33",2015,2.6,"Tirol"
"Y_GE25","AT34",2015,2.9,"Vorarlberg"
"Y_GE25","BE",2015,7.3,"Belgium"
"Y_GE25","BE1",2015,16.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2015,16.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2015,4.3,"Vlaams Gewest"
"Y_GE25","BE21",2015,5.3,"Prov. Antwerpen"
"Y_GE25","BE22",2015,5,"Prov. Limburg (BE)"
"Y_GE25","BE23",2015,3.4,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2015,4.3,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2015,3.5,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2015,10.1,"Région wallonne"
"Y_GE25","BE31",2015,6.7,"Prov. Brabant Wallon"
"Y_GE25","BE32",2015,11.2,"Prov. Hainaut"
"Y_GE25","BE33",2015,11.2,"Prov. Liège"
"Y_GE25","BE34",2015,8.3,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2015,8.8,"Prov. Namur"
"Y_GE25","BG",2015,8.4,"Bulgaria"
"Y_GE25","BG3",2015,9.9,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2015,11.1,"Severozapaden"
"Y_GE25","BG32",2015,9.9,"Severen tsentralen"
"Y_GE25","BG33",2015,9.6,"Severoiztochen"
"Y_GE25","BG34",2015,9.3,"Yugoiztochen"
"Y_GE25","BG4",2015,7.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2015,6.2,"Yugozapaden"
"Y_GE25","BG42",2015,8.4,"Yuzhen tsentralen"
"Y_GE25","CH",2015,4,"Switzerland"
"Y_GE25","CH0",2015,4,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2015,5.8,"Région lémanique"
"Y_GE25","CH02",2015,3.6,"Espace Mittelland"
"Y_GE25","CH03",2015,3.4,"Nordwestschweiz"
"Y_GE25","CH04",2015,3.7,"Zürich"
"Y_GE25","CH05",2015,3.4,"Ostschweiz"
"Y_GE25","CH06",2015,2.9,"Zentralschweiz"
"Y_GE25","CH07",2015,5.8,"Ticino"
"Y_GE25","CY",2015,13.2,"Cyprus"
"Y_GE25","CY0",2015,13.2,"Kypros"
"Y_GE25","CY00",2015,13.2,"Kypros"
"Y_GE25","CZ",2015,4.5,"Czech Republic"
"Y_GE25","CZ0",2015,4.5,"Ceská republika"
"Y_GE25","CZ01",2015,2.5,"Praha"
"Y_GE25","CZ02",2015,2.9,"Strední Cechy"
"Y_GE25","CZ03",2015,3.5,"Jihozápad"
"Y_GE25","CZ04",2015,6.5,"Severozápad"
"Y_GE25","CZ05",2015,4.7,"Severovýchod"
"Y_GE25","CZ06",2015,4.3,"Jihovýchod"
"Y_GE25","CZ07",2015,5,"Strední Morava"
"Y_GE25","CZ08",2015,7.5,"Moravskoslezsko"
"Y_GE25","DE",2015,4.3,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2015,2.7,"Baden-Württemberg"
"Y_GE25","DE11",2015,2.9,"Stuttgart"
"Y_GE25","DE12",2015,3,"Karlsruhe"
"Y_GE25","DE13",2015,2.2,"Freiburg"
"Y_GE25","DE14",2015,2.6,"Tübingen"
"Y_GE25","DE2",2015,2.7,"Bayern"
"Y_GE25","DE21",2015,2.6,"Oberbayern"
"Y_GE25","DE22",2015,2.4,"Niederbayern"
"Y_GE25","DE23",2015,2.5,"Oberpfalz"
"Y_GE25","DE24",2015,3.6,"Oberfranken"
"Y_GE25","DE25",2015,2.8,"Mittelfranken"
"Y_GE25","DE26",2015,2.7,"Unterfranken"
"Y_GE25","DE27",2015,2.8,"Schwaben"
"Y_GE25","DE3",2015,8.9,"Berlin"
"Y_GE25","DE30",2015,8.9,"Berlin"
"Y_GE25","DE4",2015,5.6,"Brandenburg"
"Y_GE25","DE40",2015,5.6,"Brandenburg"
"Y_GE25","DE5",2015,5.2,"Bremen"
"Y_GE25","DE50",2015,5.2,"Bremen"
"Y_GE25","DE6",2015,4,"Hamburg"
"Y_GE25","DE60",2015,4,"Hamburg"
"Y_GE25","DE7",2015,3.7,"Hessen"
"Y_GE25","DE71",2015,3.8,"Darmstadt"
"Y_GE25","DE72",2015,3.4,"Gießen"
"Y_GE25","DE73",2015,3.3,"Kassel"
"Y_GE25","DE8",2015,7.6,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2015,7.6,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2015,4,"Niedersachsen"
"Y_GE25","DE91",2015,4.8,"Braunschweig"
"Y_GE25","DE92",2015,4.4,"Hannover"
"Y_GE25","DE93",2015,3.2,"Lüneburg"
"Y_GE25","DE94",2015,3.7,"Weser-Ems"
"Y_GE25","DEA",2015,4.9,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2015,5.6,"Düsseldorf"
"Y_GE25","DEA2",2015,4.6,"Köln"
"Y_GE25","DEA3",2015,3.9,"Münster"
"Y_GE25","DEA4",2015,4.2,"Detmold"
"Y_GE25","DEA5",2015,5.2,"Arnsberg"
"Y_GE25","DEB",2015,3.2,"Rheinland-Pfalz"
"Y_GE25","DEB1",2015,3.2,"Koblenz"
"Y_GE25","DEB2",2015,2.5,"Trier"
"Y_GE25","DEB3",2015,3.4,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2015,5.1,"Saarland"
"Y_GE25","DEC0",2015,5.1,"Saarland"
"Y_GE25","DED",2015,6.1,"Sachsen"
"Y_GE25","DED2",2015,6,"Dresden"
"Y_GE25","DED4",2015,5.3,"Chemnitz"
"Y_GE25","DED5",2015,7.6,"Leipzig"
"Y_GE25","DEE",2015,7.7,"Sachsen-Anhalt"
"Y_GE25","DEE0",2015,7.7,"Sachsen-Anhalt"
"Y_GE25","DEF",2015,3.7,"Schleswig-Holstein"
"Y_GE25","DEF0",2015,3.7,"Schleswig-Holstein"
"Y_GE25","DEG",2015,5.5,"Thüringen"
"Y_GE25","DEG0",2015,5.5,"Thüringen"
"Y_GE25","DK",2015,5.3,"Denmark"
"Y_GE25","DK0",2015,5.3,"Danmark"
"Y_GE25","DK01",2015,6.1,"Hovedstaden"
"Y_GE25","DK02",2015,5,"Sjælland"
"Y_GE25","DK03",2015,5.1,"Syddanmark"
"Y_GE25","DK04",2015,4.7,"Midtjylland"
"Y_GE25","DK05",2015,5.1,"Nordjylland"
"Y_GE25","EA17",2015,9.7,"Euro area (17 countries)"
"Y_GE25","EA18",2015,9.7,"Euro area (18 countries)"
"Y_GE25","EA19",2015,9.7,"Euro area (19 countries)"
"Y_GE25","EE",2015,5.6,"Estonia"
"Y_GE25","EE0",2015,5.6,"Eesti"
"Y_GE25","EE00",2015,5.6,"Eesti"
"Y_GE25","EL",2015,23.4,"Greece"
"Y_GE25","EL3",2015,23.9,"Attiki"
"Y_GE25","EL30",2015,23.9,"Attiki"
"Y_GE25","EL4",2015,19.1,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2015,16.1,"Voreio Aigaio"
"Y_GE25","EL42",2015,13.3,"Notio Aigaio"
"Y_GE25","EL43",2015,23.2,"Kriti"
"Y_GE25","EL5",2015,24.1,"Voreia Ellada"
"Y_GE25","EL51",2015,21,"Anatoliki Makedonia, Thraki"
"Y_GE25","EL52",2015,24.6,"Kentriki Makedonia"
"Y_GE25","EL53",2015,29.3,"Dytiki Makedonia"
"Y_GE25","EL54",2015,23,"Ipeiros"
"Y_GE25","EL6",2015,23.4,"Kentriki Ellada"
"Y_GE25","EL61",2015,24.7,"Thessalia"
"Y_GE25","EL62",2015,16.6,"Ionia Nisia"
"Y_GE25","EL63",2015,26.4,"Dytiki Ellada"
"Y_GE25","EL64",2015,23.6,"Sterea Ellada"
"Y_GE25","EL65",2015,20.8,"Peloponnisos"
"Y_GE25","ES",2015,20.1,"Spain"
"Y_GE25","ES1",2015,17.8,"Noroeste (ES)"
"Y_GE25","ES11",2015,18,"Galicia"
"Y_GE25","ES12",2015,18.1,"Principado de Asturias"
"Y_GE25","ES13",2015,16.6,"Cantabria"
"Y_GE25","ES2",2015,13.7,"Noreste (ES)"
"Y_GE25","ES21",2015,13.5,"País Vasco"
"Y_GE25","ES22",2015,12.4,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2015,13.9,"La Rioja"
"Y_GE25","ES24",2015,14.7,"Aragón"
"Y_GE25","ES3",2015,15.2,"Comunidad de Madrid"
"Y_GE25","ES30",2015,15.2,"Comunidad de Madrid"
"Y_GE25","ES4",2015,21.2,"Centro (ES)"
"Y_GE25","ES41",2015,16.6,"Castilla y León"
"Y_GE25","ES42",2015,23.8,"Castilla-la Mancha"
"Y_GE25","ES43",2015,26.9,"Extremadura"
"Y_GE25","ES5",2015,18.1,"Este (ES)"
"Y_GE25","ES51",2015,16.8,"Cataluña"
"Y_GE25","ES52",2015,20.8,"Comunidad Valenciana"
"Y_GE25","ES53",2015,15.4,"Illes Balears"
"Y_GE25","ES6",2015,28.3,"Sur (ES)"
"Y_GE25","ES61",2015,29.4,"Andalucía"
"Y_GE25","ES62",2015,22.3,"Región de Murcia"
"Y_GE25","ES63",2015,22.4,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2015,29.8,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2015,27.3,"Canarias (ES)"
"Y_GE25","ES70",2015,27.3,"Canarias (ES)"
"Y_GE25","EU15",2015,8.6,"European Union (15 countries)"
"Y_GE25","EU27",2015,8.2,"European Union (27 countries)"
"Y_GE25","EU28",2015,8.3,"European Union (28 countries)"
"Y_GE25","FI",2015,7.6,"Finland"
"Y_GE25","FI1",2015,7.6,"Manner-Suomi"
"Y_GE25","FI19",2015,7.7,"Länsi-Suomi"
"Y_GE25","FI1B",2015,6.6,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2015,8.3,"Etelä-Suomi"
"Y_GE25","FI1D",2015,8.3,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2015,NA,"Åland"
"Y_GE25","FI20",2015,NA,"Åland"
"Y_GE25","FR",2015,8.9,"France"
"Y_GE25","FR1",2015,8.3,"Île de France"
"Y_GE25","FR10",2015,8.3,"Île de France"
"Y_GE25","FR2",2015,8.8,"Bassin Parisien"
"Y_GE25","FR21",2015,10.9,"Champagne-Ardenne"
"Y_GE25","FR22",2015,9.2,"Picardie"
"Y_GE25","FR23",2015,9,"Haute-Normandie"
"Y_GE25","FR24",2015,9.3,"Centre (FR)"
"Y_GE25","FR25",2015,7.1,"Basse-Normandie"
"Y_GE25","FR26",2015,7,"Bourgogne"
"Y_GE25","FR3",2015,12.1,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2015,12.1,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2015,8.5,"Est (FR)"
"Y_GE25","FR41",2015,10.1,"Lorraine"
"Y_GE25","FR42",2015,7.3,"Alsace"
"Y_GE25","FR43",2015,7.3,"Franche-Comté"
"Y_GE25","FR5",2015,7.3,"Ouest (FR)"
"Y_GE25","FR51",2015,7.4,"Pays de la Loire"
"Y_GE25","FR52",2015,6.7,"Bretagne"
"Y_GE25","FR53",2015,8.2,"Poitou-Charentes"
"Y_GE25","FR6",2015,7.8,"Sud-Ouest (FR)"
"Y_GE25","FR61",2015,8.3,"Aquitaine"
"Y_GE25","FR62",2015,7.3,"Midi-Pyrénées"
"Y_GE25","FR63",2015,7.3,"Limousin"
"Y_GE25","FR7",2015,7.8,"Centre-Est (FR)"
"Y_GE25","FR71",2015,7.8,"Rhône-Alpes"
"Y_GE25","FR72",2015,7.6,"Auvergne"
"Y_GE25","FR8",2015,10.2,"Méditerranée"
"Y_GE25","FR81",2015,11.1,"Languedoc-Roussillon"
"Y_GE25","FR82",2015,9.8,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2015,NA,"Corse"
"Y_GE25","FRA",2015,19.7,"Départements d'outre-mer"
"Y_GE25","FRA1",2015,21.3,"Guadeloupe"
"Y_GE25","FRA2",2015,16.7,"Martinique"
"Y_GE25","FRA3",2015,18.9,"Guyane"
"Y_GE25","FRA4",2015,20.6,"La Réunion"
"Y_GE25","FRA5",2015,20,"Mayotte"
"Y_GE25","HR",2015,13.8,"Croatia"
"Y_GE25","HR0",2015,13.8,"Hrvatska"
"Y_GE25","HR03",2015,14.4,"Jadranska Hrvatska"
"Y_GE25","HR04",2015,13.5,"Kontinentalna Hrvatska"
"Y_GE25","HU",2015,6,"Hungary"
"Y_GE25","HU1",2015,4.9,"Közép-Magyarország"
"Y_GE25","HU10",2015,4.9,"Közép-Magyarország"
"Y_GE25","HU2",2015,4.6,"Dunántúl"
"Y_GE25","HU21",2015,4,"Közép-Dunántúl"
"Y_GE25","HU22",2015,3.1,"Nyugat-Dunántúl"
"Y_GE25","HU23",2015,7.2,"Dél-Dunántúl"
"Y_GE25","HU3",2015,8,"Alföld és Észak"
"Y_GE25","HU31",2015,7.6,"Észak-Magyarország"
"Y_GE25","HU32",2015,9.5,"Észak-Alföld"
"Y_GE25","HU33",2015,6.7,"Dél-Alföld"
"Y_GE25","IE",2015,8.3,"Ireland"
"Y_GE25","IE0",2015,8.3,"Éire/Ireland"
"Y_GE25","IE01",2015,9.2,"Border, Midland and Western"
"Y_GE25","IE02",2015,8,"Southern and Eastern"
"Y_GE25","IS",2015,3,"Iceland"
"Y_GE25","IS0",2015,3,"Ísland"
"Y_GE25","IS00",2015,3,"Ísland"
"Y_GE25","IT",2015,10.1,"Italy"
"Y_GE25","ITC",2015,7.1,"Nord-Ovest"
"Y_GE25","ITC1",2015,8.5,"Piemonte"
"Y_GE25","ITC2",2015,7.4,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2015,8,"Liguria"
"Y_GE25","ITC4",2015,6.4,"Lombardia"
"Y_GE25","ITF",2015,16.2,"Sud"
"Y_GE25","ITF1",2015,10.4,"Abruzzo"
"Y_GE25","ITF2",2015,12.7,"Molise"
"Y_GE25","ITF3",2015,17,"Campania"
"Y_GE25","ITF4",2015,16.9,"Puglia"
"Y_GE25","ITF5",2015,11.3,"Basilicata"
"Y_GE25","ITF6",2015,19.6,"Calabria"
"Y_GE25","ITG",2015,17.3,"Isole"
"Y_GE25","ITG1",2015,18.3,"Sicilia"
"Y_GE25","ITG2",2015,14.8,"Sardegna"
"Y_GE25","ITH",2015,6.2,"Nord-Est"
"Y_GE25","ITH1",2015,3.1,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2015,5.7,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2015,6,"Veneto"
"Y_GE25","ITH4",2015,6.9,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2015,6.5,"Emilia-Romagna"
"Y_GE25","ITI",2015,9.1,"Centro (IT)"
"Y_GE25","ITI1",2015,7.9,"Toscana"
"Y_GE25","ITI2",2015,8.7,"Umbria"
"Y_GE25","ITI3",2015,8.6,"Marche"
"Y_GE25","ITI4",2015,10.2,"Lazio"
"Y_GE25","LT",2015,8.5,"Lithuania"
"Y_GE25","LT0",2015,8.5,"Lietuva"
"Y_GE25","LT00",2015,8.5,"Lietuva"
"Y_GE25","LU",2015,5.7,"Luxembourg"
"Y_GE25","LU0",2015,5.7,"Luxembourg"
"Y_GE25","LU00",2015,5.7,"Luxembourg"
"Y_GE25","LV",2015,9.3,"Latvia"
"Y_GE25","LV0",2015,9.3,"Latvija"
"Y_GE25","LV00",2015,9.3,"Latvija"
"Y_GE25","MK",2015,23.8,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2015,23.8,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2015,23.8,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2015,4.4,"Malta"
"Y_GE25","MT0",2015,4.4,"Malta"
"Y_GE25","MT00",2015,4.4,"Malta"
"Y_GE25","NL",2015,6.1,"Netherlands"
"Y_GE25","NL1",2015,7.1,"Noord-Nederland"
"Y_GE25","NL11",2015,8.2,"Groningen"
"Y_GE25","NL12",2015,6.6,"Friesland (NL)"
"Y_GE25","NL13",2015,6.6,"Drenthe"
"Y_GE25","NL2",2015,5.8,"Oost-Nederland"
"Y_GE25","NL21",2015,6,"Overijssel"
"Y_GE25","NL22",2015,5.6,"Gelderland"
"Y_GE25","NL23",2015,6.7,"Flevoland"
"Y_GE25","NL3",2015,6.1,"West-Nederland"
"Y_GE25","NL31",2015,5.5,"Utrecht"
"Y_GE25","NL32",2015,5.7,"Noord-Holland"
"Y_GE25","NL33",2015,6.8,"Zuid-Holland"
"Y_GE25","NL34",2015,4.8,"Zeeland"
"Y_GE25","NL4",2015,5.7,"Zuid-Nederland"
"Y_GE25","NL41",2015,5.7,"Noord-Brabant"
"Y_GE25","NL42",2015,5.5,"Limburg (NL)"
"Y_GE25","NO",2015,3.4,"Norway"
"Y_GE25","NO0",2015,3.4,"Norge"
"Y_GE25","NO01",2015,4.1,"Oslo og Akershus"
"Y_GE25","NO02",2015,3.8,"Hedmark og Oppland"
"Y_GE25","NO03",2015,3.4,"Sør-Østlandet"
"Y_GE25","NO04",2015,3.9,"Agder og Rogaland"
"Y_GE25","NO05",2015,3,"Vestlandet"
"Y_GE25","NO06",2015,2.7,"Trøndelag"
"Y_GE25","NO07",2015,2,"Nord-Norge"
"Y_GE25","PL",2015,6.4,"Poland"
"Y_GE25","PL1",2015,5.9,"Region Centralny"
"Y_GE25","PL11",2015,6.6,"Lódzkie"
"Y_GE25","PL12",2015,5.5,"Mazowieckie"
"Y_GE25","PL2",2015,6.1,"Region Poludniowy"
"Y_GE25","PL21",2015,5.8,"Malopolskie"
"Y_GE25","PL22",2015,6.3,"Slaskie"
"Y_GE25","PL3",2015,8.1,"Region Wschodni"
"Y_GE25","PL31",2015,7.9,"Lubelskie"
"Y_GE25","PL32",2015,9.3,"Podkarpackie"
"Y_GE25","PL33",2015,8.4,"Swietokrzyskie"
"Y_GE25","PL34",2015,6,"Podlaskie"
"Y_GE25","PL4",2015,5.3,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2015,4.7,"Wielkopolskie"
"Y_GE25","PL42",2015,6.3,"Zachodniopomorskie"
"Y_GE25","PL43",2015,5.7,"Lubuskie"
"Y_GE25","PL5",2015,6,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2015,6.2,"Dolnoslaskie"
"Y_GE25","PL52",2015,5.7,"Opolskie"
"Y_GE25","PL6",2015,6.6,"Region Pólnocny"
"Y_GE25","PL61",2015,6.8,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2015,8.3,"Warminsko-Mazurskie"
"Y_GE25","PL63",2015,5.4,"Pomorskie"
"Y_GE25","PT",2015,11,"Portugal"
"Y_GE25","PT1",2015,10.9,"Continente"
"Y_GE25","PT11",2015,12,"Norte"
"Y_GE25","PT15",2015,11.2,"Algarve"
"Y_GE25","PT16",2015,7.9,"Centro (PT)"
"Y_GE25","PT17",2015,11.8,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2015,11.7,"Alentejo"
"Y_GE25","PT2",2015,10.5,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2015,10.5,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2015,12.4,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2015,12.4,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2015,5.6,"Romania"
"Y_GE25","RO1",2015,4.6,"Macroregiunea unu"
"Y_GE25","RO11",2015,3.7,"Nord-Vest"
"Y_GE25","RO12",2015,5.9,"Centru"
"Y_GE25","RO2",2015,4.7,"Macroregiunea doi"
"Y_GE25","RO21",2015,3,"Nord-Est"
"Y_GE25","RO22",2015,7.3,"Sud-Est"
"Y_GE25","RO3",2015,6.7,"Macroregiunea trei"
"Y_GE25","RO31",2015,8.3,"Sud - Muntenia"
"Y_GE25","RO32",2015,4.8,"Bucuresti - Ilfov"
"Y_GE25","RO4",2015,6.7,"Macroregiunea patru"
"Y_GE25","RO41",2015,8.7,"Sud-Vest Oltenia"
"Y_GE25","RO42",2015,4.3,"Vest"
"Y_GE25","SE",2015,5.6,"Sweden"
"Y_GE25","SE1",2015,5.6,"Östra Sverige"
"Y_GE25","SE11",2015,5.5,"Stockholm"
"Y_GE25","SE12",2015,5.7,"Östra Mellansverige"
"Y_GE25","SE2",2015,5.6,"Södra Sverige"
"Y_GE25","SE21",2015,4.1,"Småland med öarna"
"Y_GE25","SE22",2015,7.6,"Sydsverige"
"Y_GE25","SE23",2015,4.8,"Västsverige"
"Y_GE25","SE3",2015,5.4,"Norra Sverige"
"Y_GE25","SE31",2015,5.7,"Norra Mellansverige"
"Y_GE25","SE32",2015,5.2,"Mellersta Norrland"
"Y_GE25","SE33",2015,5.2,"Övre Norrland"
"Y_GE25","SI",2015,8.4,"Slovenia"
"Y_GE25","SI0",2015,8.4,"Slovenija"
"Y_GE25","SI03",2015,9.8,"Vzhodna Slovenija"
"Y_GE25","SI04",2015,6.8,"Zahodna Slovenija"
"Y_GE25","SK",2015,10.2,"Slovakia"
"Y_GE25","SK0",2015,10.2,"Slovensko"
"Y_GE25","SK01",2015,5.2,"Bratislavský kraj"
"Y_GE25","SK02",2015,8.8,"Západné Slovensko"
"Y_GE25","SK03",2015,11.2,"Stredné Slovensko"
"Y_GE25","SK04",2015,13.5,"Východné Slovensko"
"Y_GE25","TR",2015,8.6,"Turkey"
"Y_GE25","TR1",2015,11.3,"Istanbul"
"Y_GE25","TR10",2015,11.3,"Istanbul"
"Y_GE25","TR2",2015,5.3,"Bati Marmara"
"Y_GE25","TR21",2015,6.1,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2015,4.4,"Balikesir, Çanakkale"
"Y_GE25","TR3",2015,8,"Ege"
"Y_GE25","TR31",2015,13.2,"Izmir"
"Y_GE25","TR32",2015,5.6,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2015,3.1,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2015,7.3,"Dogu Marmara"
"Y_GE25","TR41",2015,6.3,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2015,8.2,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2015,8.3,"Bati Anadolu"
"Y_GE25","TR51",2015,9.5,"Ankara"
"Y_GE25","TR52",2015,5.1,"Konya, Karaman"
"Y_GE25","TR6",2015,9.5,"Akdeniz"
"Y_GE25","TR61",2015,8.1,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2015,8.4,"Adana, Mersin"
"Y_GE25","TR63",2015,13.3,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2015,7.8,"Orta Anadolu"
"Y_GE25","TR71",2015,7.8,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2015,7.8,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2015,5.4,"Bati Karadeniz"
"Y_GE25","TR81",2015,5.3,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2015,5.4,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2015,5.5,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2015,3.5,"Dogu Karadeniz"
"Y_GE25","TR90",2015,3.5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2015,4.1,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2015,5.1,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2015,3.1,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2015,7.4,"Ortadogu Anadolu"
"Y_GE25","TRB1",2015,6,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2015,9,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2015,14,"Güneydogu Anadolu"
"Y_GE25","TRC1",2015,8,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2015,16.3,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2015,20,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2015,3.8,"United Kingdom"
"Y_GE25","UKC",2015,5.8,"North East (UK)"
"Y_GE25","UKC1",2015,5.8,"Tees Valley and Durham"
"Y_GE25","UKC2",2015,5.8,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2015,4,"North West (UK)"
"Y_GE25","UKD1",2015,3.4,"Cumbria"
"Y_GE25","UKD3",2015,4.8,"Greater Manchester"
"Y_GE25","UKD4",2015,3.6,"Lancashire"
"Y_GE25","UKD6",2015,2.5,"Cheshire"
"Y_GE25","UKD7",2015,4.3,"Merseyside"
"Y_GE25","UKE",2015,4.4,"Yorkshire and The Humber"
"Y_GE25","UKE1",2015,4.9,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2015,1.6,"North Yorkshire"
"Y_GE25","UKE3",2015,5.9,"South Yorkshire"
"Y_GE25","UKE4",2015,4.5,"West Yorkshire"
"Y_GE25","UKF",2015,3.5,"East Midlands (UK)"
"Y_GE25","UKF1",2015,3.8,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2015,3.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2015,3,"Lincolnshire"
"Y_GE25","UKG",2015,4.3,"West Midlands (UK)"
"Y_GE25","UKG1",2015,2.3,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2015,3.5,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2015,6,"West Midlands"
"Y_GE25","UKH",2015,3,"East of England"
"Y_GE25","UKH1",2015,3.1,"East Anglia"
"Y_GE25","UKH2",2015,2.7,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2015,3.2,"Essex"
"Y_GE25","UKI",2015,4.7,"London"
"Y_GE25","UKI3",2015,4.6,"Inner London - West"
"Y_GE25","UKI4",2015,5.3,"Inner London - East"
"Y_GE25","UKI5",2015,5.4,"Outer London - East and North East"
"Y_GE25","UKI6",2015,3.5,"Outer London - South"
"Y_GE25","UKI7",2015,4,"Outer London - West and North West"
"Y_GE25","UKJ",2015,2.8,"South East (UK)"
"Y_GE25","UKJ1",2015,2.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2015,2.4,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2015,2.8,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2015,3.7,"Kent"
"Y_GE25","UKK",2015,2.7,"South West (UK)"
"Y_GE25","UKK1",2015,2.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2015,2.5,"Dorset and Somerset"
"Y_GE25","UKK3",2015,2.8,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2015,2.4,"Devon"
"Y_GE25","UKL",2015,3.6,"Wales"
"Y_GE25","UKL1",2015,4.1,"West Wales and The Valleys"
"Y_GE25","UKL2",2015,2.8,"East Wales"
"Y_GE25","UKM",2015,4.2,"Scotland"
"Y_GE25","UKM2",2015,4.1,"Eastern Scotland"
"Y_GE25","UKM3",2015,5.1,"South Western Scotland"
"Y_GE25","UKM5",2015,2.2,"North Eastern Scotland"
"Y_GE25","UKM6",2015,3.4,"Highlands and Islands"
"Y_GE25","UKN",2015,4.1,"Northern Ireland (UK)"
"Y_GE25","UKN0",2015,4.1,"Northern Ireland (UK)"
"Y15-24","AT",2014,10.3,"Austria"
"Y15-24","AT1",2014,14.2,"Ostösterreich"
"Y15-24","AT11",2014,NA,"Burgenland (AT)"
"Y15-24","AT12",2014,11.1,"Niederösterreich"
"Y15-24","AT13",2014,18,"Wien"
"Y15-24","AT2",2014,8.4,"Südösterreich"
"Y15-24","AT21",2014,9.4,"Kärnten"
"Y15-24","AT22",2014,7.9,"Steiermark"
"Y15-24","AT3",2014,7.3,"Westösterreich"
"Y15-24","AT31",2014,7.9,"Oberösterreich"
"Y15-24","AT32",2014,NA,"Salzburg"
"Y15-24","AT33",2014,6,"Tirol"
"Y15-24","AT34",2014,NA,"Vorarlberg"
"Y15-24","BE",2014,23.2,"Belgium"
"Y15-24","BE1",2014,39.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2014,39.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2014,16.1,"Vlaams Gewest"
"Y15-24","BE21",2014,17.9,"Prov. Antwerpen"
"Y15-24","BE22",2014,14.7,"Prov. Limburg (BE)"
"Y15-24","BE23",2014,16,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2014,18.5,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2014,13.2,"Prov. West-Vlaanderen"
"Y15-24","BE3",2014,32.1,"Région wallonne"
"Y15-24","BE31",2014,25.1,"Prov. Brabant Wallon"
"Y15-24","BE32",2014,36.7,"Prov. Hainaut"
"Y15-24","BE33",2014,32.3,"Prov. Liège"
"Y15-24","BE34",2014,23.2,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2014,29.9,"Prov. Namur"
"Y15-24","BG",2014,23.8,"Bulgaria"
"Y15-24","BG3",2014,25.8,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2014,27.7,"Severozapaden"
"Y15-24","BG32",2014,24.9,"Severen tsentralen"
"Y15-24","BG33",2014,22.6,"Severoiztochen"
"Y15-24","BG34",2014,28.6,"Yugoiztochen"
"Y15-24","BG4",2014,21.8,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2014,16.8,"Yugozapaden"
"Y15-24","BG42",2014,28.9,"Yuzhen tsentralen"
"Y15-24","CH",2014,8.6,"Switzerland"
"Y15-24","CH0",2014,8.6,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2014,14.3,"Région lémanique"
"Y15-24","CH02",2014,8.6,"Espace Mittelland"
"Y15-24","CH03",2014,6.5,"Nordwestschweiz"
"Y15-24","CH04",2014,6.6,"Zürich"
"Y15-24","CH05",2014,5.5,"Ostschweiz"
"Y15-24","CH06",2014,7.4,"Zentralschweiz"
"Y15-24","CH07",2014,17,"Ticino"
"Y15-24","CY",2014,36,"Cyprus"
"Y15-24","CY0",2014,36,"Kypros"
"Y15-24","CY00",2014,36,"Kypros"
"Y15-24","CZ",2014,15.9,"Czech Republic"
"Y15-24","CZ0",2014,15.9,"Ceská republika"
"Y15-24","CZ01",2014,10.1,"Praha"
"Y15-24","CZ02",2014,13.2,"Strední Cechy"
"Y15-24","CZ03",2014,15.3,"Jihozápad"
"Y15-24","CZ04",2014,22.9,"Severozápad"
"Y15-24","CZ05",2014,16.2,"Severovýchod"
"Y15-24","CZ06",2014,14.6,"Jihovýchod"
"Y15-24","CZ07",2014,14.4,"Strední Morava"
"Y15-24","CZ08",2014,18.9,"Moravskoslezsko"
"Y15-24","DE",2014,7.7,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2014,5,"Baden-Württemberg"
"Y15-24","DE11",2014,4.7,"Stuttgart"
"Y15-24","DE12",2014,4.8,"Karlsruhe"
"Y15-24","DE13",2014,5,"Freiburg"
"Y15-24","DE14",2014,5.8,"Tübingen"
"Y15-24","DE2",2014,4.4,"Bayern"
"Y15-24","DE21",2014,3.7,"Oberbayern"
"Y15-24","DE22",2014,NA,"Niederbayern"
"Y15-24","DE23",2014,NA,"Oberpfalz"
"Y15-24","DE24",2014,NA,"Oberfranken"
"Y15-24","DE25",2014,6,"Mittelfranken"
"Y15-24","DE26",2014,NA,"Unterfranken"
"Y15-24","DE27",2014,NA,"Schwaben"
"Y15-24","DE3",2014,15.5,"Berlin"
"Y15-24","DE30",2014,15.5,"Berlin"
"Y15-24","DE4",2014,10.8,"Brandenburg"
"Y15-24","DE40",2014,10.8,"Brandenburg"
"Y15-24","DE5",2014,NA,"Bremen"
"Y15-24","DE50",2014,NA,"Bremen"
"Y15-24","DE6",2014,7.8,"Hamburg"
"Y15-24","DE60",2014,7.8,"Hamburg"
"Y15-24","DE7",2014,9.5,"Hessen"
"Y15-24","DE71",2014,9.4,"Darmstadt"
"Y15-24","DE72",2014,10.7,"Gießen"
"Y15-24","DE73",2014,8.5,"Kassel"
"Y15-24","DE8",2014,11.5,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2014,11.5,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2014,6.9,"Niedersachsen"
"Y15-24","DE91",2014,7.4,"Braunschweig"
"Y15-24","DE92",2014,7.4,"Hannover"
"Y15-24","DE93",2014,6.5,"Lüneburg"
"Y15-24","DE94",2014,6.6,"Weser-Ems"
"Y15-24","DEA",2014,9.3,"Nordrhein-Westfalen"
"Y15-24","DEA1",2014,8.7,"Düsseldorf"
"Y15-24","DEA2",2014,9.6,"Köln"
"Y15-24","DEA3",2014,9.1,"Münster"
"Y15-24","DEA4",2014,9.4,"Detmold"
"Y15-24","DEA5",2014,10.1,"Arnsberg"
"Y15-24","DEB",2014,7.6,"Rheinland-Pfalz"
"Y15-24","DEB1",2014,8.1,"Koblenz"
"Y15-24","DEB2",2014,NA,"Trier"
"Y15-24","DEB3",2014,7.6,"Rheinhessen-Pfalz"
"Y15-24","DEC",2014,NA,"Saarland"
"Y15-24","DEC0",2014,NA,"Saarland"
"Y15-24","DED",2014,10.9,"Sachsen"
"Y15-24","DED2",2014,13,"Dresden"
"Y15-24","DED4",2014,NA,"Chemnitz"
"Y15-24","DED5",2014,NA,"Leipzig"
"Y15-24","DEE",2014,12.1,"Sachsen-Anhalt"
"Y15-24","DEE0",2014,12.1,"Sachsen-Anhalt"
"Y15-24","DEF",2014,8.5,"Schleswig-Holstein"
"Y15-24","DEF0",2014,8.5,"Schleswig-Holstein"
"Y15-24","DEG",2014,8.4,"Thüringen"
"Y15-24","DEG0",2014,8.4,"Thüringen"
"Y15-24","DK",2014,12.6,"Denmark"
"Y15-24","DK0",2014,12.6,"Danmark"
"Y15-24","DK01",2014,12.8,"Hovedstaden"
"Y15-24","DK02",2014,14.3,"Sjælland"
"Y15-24","DK03",2014,12.5,"Syddanmark"
"Y15-24","DK04",2014,11.5,"Midtjylland"
"Y15-24","DK05",2014,12.9,"Nordjylland"
"Y15-24","EA17",2014,23.8,"Euro area (17 countries)"
"Y15-24","EA18",2014,23.8,"Euro area (18 countries)"
"Y15-24","EA19",2014,23.8,"Euro area (19 countries)"
"Y15-24","EE",2014,15,"Estonia"
"Y15-24","EE0",2014,15,"Eesti"
"Y15-24","EE00",2014,15,"Eesti"
"Y15-24","EL",2014,52.4,"Greece"
"Y15-24","EL3",2014,52.5,"Attiki"
"Y15-24","EL30",2014,52.5,"Attiki"
"Y15-24","EL4",2014,38.9,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2014,40.2,"Voreio Aigaio"
"Y15-24","EL42",2014,25.8,"Notio Aigaio"
"Y15-24","EL43",2014,46.3,"Kriti"
"Y15-24","EL5",2014,54.1,"Voreia Ellada"
"Y15-24","EL51",2014,50.7,"Anatoliki Makedonia, Thraki"
"Y15-24","EL52",2014,53.4,"Kentriki Makedonia"
"Y15-24","EL53",2014,49.6,"Dytiki Makedonia"
"Y15-24","EL54",2014,69.8,"Ipeiros"
"Y15-24","EL6",2014,57.3,"Kentriki Ellada"
"Y15-24","EL61",2014,59.8,"Thessalia"
"Y15-24","EL62",2014,44.8,"Ionia Nisia"
"Y15-24","EL63",2014,61.1,"Dytiki Ellada"
"Y15-24","EL64",2014,59.1,"Sterea Ellada"
"Y15-24","EL65",2014,52,"Peloponnisos"
"Y15-24","ES",2014,53.2,"Spain"
"Y15-24","ES1",2014,47.8,"Noroeste (ES)"
"Y15-24","ES11",2014,48.5,"Galicia"
"Y15-24","ES12",2014,45.1,"Principado de Asturias"
"Y15-24","ES13",2014,49.2,"Cantabria"
"Y15-24","ES2",2014,47.3,"Noreste (ES)"
"Y15-24","ES21",2014,45,"País Vasco"
"Y15-24","ES22",2014,45.2,"Comunidad Foral de Navarra"
"Y15-24","ES23",2014,44.8,"La Rioja"
"Y15-24","ES24",2014,51.5,"Aragón"
"Y15-24","ES3",2014,49,"Comunidad de Madrid"
"Y15-24","ES30",2014,49,"Comunidad de Madrid"
"Y15-24","ES4",2014,56.3,"Centro (ES)"
"Y15-24","ES41",2014,50.4,"Castilla y León"
"Y15-24","ES42",2014,61.3,"Castilla-la Mancha"
"Y15-24","ES43",2014,55.4,"Extremadura"
"Y15-24","ES5",2014,50.2,"Este (ES)"
"Y15-24","ES51",2014,47.1,"Cataluña"
"Y15-24","ES52",2014,56.7,"Comunidad Valenciana"
"Y15-24","ES53",2014,44.4,"Illes Balears"
"Y15-24","ES6",2014,60.2,"Sur (ES)"
"Y15-24","ES61",2014,61.5,"Andalucía"
"Y15-24","ES62",2014,52.4,"Región de Murcia"
"Y15-24","ES63",2014,67.5,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2014,57.3,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2014,57.4,"Canarias (ES)"
"Y15-24","ES70",2014,57.4,"Canarias (ES)"
"Y15-24","EU15",2014,21.9,"European Union (15 countries)"
"Y15-24","EU27",2014,22,"European Union (27 countries)"
"Y15-24","EU28",2014,22.2,"European Union (28 countries)"
"Y15-24","FI",2014,20.5,"Finland"
"Y15-24","FI1",2014,20.6,"Manner-Suomi"
"Y15-24","FI19",2014,20.1,"Länsi-Suomi"
"Y15-24","FI1B",2014,18.3,"Helsinki-Uusimaa"
"Y15-24","FI1C",2014,22.9,"Etelä-Suomi"
"Y15-24","FI1D",2014,22.1,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2014,NA,"Åland"
"Y15-24","FI20",2014,NA,"Åland"
"Y15-24","FR",2014,24.3,"France"
"Y15-24","FR1",2014,21.4,"Île de France"
"Y15-24","FR10",2014,21.4,"Île de France"
"Y15-24","FR2",2014,24.1,"Bassin Parisien"
"Y15-24","FR21",2014,25.2,"Champagne-Ardenne"
"Y15-24","FR22",2014,27.4,"Picardie"
"Y15-24","FR23",2014,25.7,"Haute-Normandie"
"Y15-24","FR24",2014,21.4,"Centre (FR)"
"Y15-24","FR25",2014,21.2,"Basse-Normandie"
"Y15-24","FR26",2014,24,"Bourgogne"
"Y15-24","FR3",2014,29.2,"Nord - Pas-de-Calais"
"Y15-24","FR30",2014,29.2,"Nord - Pas-de-Calais"
"Y15-24","FR4",2014,24.6,"Est (FR)"
"Y15-24","FR41",2014,25.7,"Lorraine"
"Y15-24","FR42",2014,25.3,"Alsace"
"Y15-24","FR43",2014,20.6,"Franche-Comté"
"Y15-24","FR5",2014,22.1,"Ouest (FR)"
"Y15-24","FR51",2014,21.3,"Pays de la Loire"
"Y15-24","FR52",2014,20.3,"Bretagne"
"Y15-24","FR53",2014,25.9,"Poitou-Charentes"
"Y15-24","FR6",2014,23.6,"Sud-Ouest (FR)"
"Y15-24","FR61",2014,23.9,"Aquitaine"
"Y15-24","FR62",2014,22.7,"Midi-Pyrénées"
"Y15-24","FR63",2014,25.2,"Limousin"
"Y15-24","FR7",2014,19.8,"Centre-Est (FR)"
"Y15-24","FR71",2014,19.8,"Rhône-Alpes"
"Y15-24","FR72",2014,20,"Auvergne"
"Y15-24","FR8",2014,27.2,"Méditerranée"
"Y15-24","FR81",2014,31.2,"Languedoc-Roussillon"
"Y15-24","FR82",2014,25.2,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2014,NA,"Corse"
"Y15-24","FRA",2014,52.2,"Départements d'outre-mer"
"Y15-24","FRA1",2014,57.3,"Guadeloupe"
"Y15-24","FRA2",2014,51.4,"Martinique"
"Y15-24","FRA3",2014,39.6,"Guyane"
"Y15-24","FRA4",2014,53.7,"La Réunion"
"Y15-24","FRA5",2014,NA,"Mayotte"
"Y15-24","HR",2014,45.5,"Croatia"
"Y15-24","HR0",2014,45.5,"Hrvatska"
"Y15-24","HR03",2014,46.5,"Jadranska Hrvatska"
"Y15-24","HR04",2014,45,"Kontinentalna Hrvatska"
"Y15-24","HU",2014,20.4,"Hungary"
"Y15-24","HU1",2014,16.1,"Közép-Magyarország"
"Y15-24","HU10",2014,16.1,"Közép-Magyarország"
"Y15-24","HU2",2014,15.3,"Dunántúl"
"Y15-24","HU21",2014,15.4,"Közép-Dunántúl"
"Y15-24","HU22",2014,12.8,"Nyugat-Dunántúl"
"Y15-24","HU23",2014,18.1,"Dél-Dunántúl"
"Y15-24","HU3",2014,26.5,"Alföld és Észak"
"Y15-24","HU31",2014,25.6,"Észak-Magyarország"
"Y15-24","HU32",2014,28.9,"Észak-Alföld"
"Y15-24","HU33",2014,24.2,"Dél-Alföld"
"Y15-24","IE",2014,23.9,"Ireland"
"Y15-24","IE0",2014,23.9,"Éire/Ireland"
"Y15-24","IE01",2014,28.7,"Border, Midland and Western"
"Y15-24","IE02",2014,22.3,"Southern and Eastern"
"Y15-24","IS",2014,9.8,"Iceland"
"Y15-24","IS0",2014,9.8,"Ísland"
"Y15-24","IS00",2014,9.8,"Ísland"
"Y15-24","IT",2014,42.7,"Italy"
"Y15-24","ITC",2014,35.5,"Nord-Ovest"
"Y15-24","ITC1",2014,42.2,"Piemonte"
"Y15-24","ITC2",2014,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2014,45,"Liguria"
"Y15-24","ITC4",2014,31.2,"Lombardia"
"Y15-24","ITF",2014,56.1,"Sud"
"Y15-24","ITF1",2014,47.4,"Abruzzo"
"Y15-24","ITF2",2014,49.3,"Molise"
"Y15-24","ITF3",2014,56,"Campania"
"Y15-24","ITF4",2014,58.1,"Puglia"
"Y15-24","ITF5",2014,46.6,"Basilicata"
"Y15-24","ITF6",2014,59.7,"Calabria"
"Y15-24","ITG",2014,55.3,"Isole"
"Y15-24","ITG1",2014,57,"Sicilia"
"Y15-24","ITG2",2014,50,"Sardegna"
"Y15-24","ITH",2014,29,"Nord-Est"
"Y15-24","ITH1",2014,12.4,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2014,27.1,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2014,27.6,"Veneto"
"Y15-24","ITH4",2014,27.1,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2014,34.9,"Emilia-Romagna"
"Y15-24","ITI",2014,42.4,"Centro (IT)"
"Y15-24","ITI1",2014,35.7,"Toscana"
"Y15-24","ITI2",2014,42.5,"Umbria"
"Y15-24","ITI3",2014,36.4,"Marche"
"Y15-24","ITI4",2014,49,"Lazio"
"Y15-24","LT",2014,19.3,"Lithuania"
"Y15-24","LT0",2014,19.3,"Lietuva"
"Y15-24","LT00",2014,19.3,"Lietuva"
"Y15-24","LU",2014,22.6,"Luxembourg"
"Y15-24","LU0",2014,22.6,"Luxembourg"
"Y15-24","LU00",2014,22.6,"Luxembourg"
"Y15-24","LV",2014,19.6,"Latvia"
"Y15-24","LV0",2014,19.6,"Latvija"
"Y15-24","LV00",2014,19.6,"Latvija"
"Y15-24","MK",2014,53.1,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2014,53.1,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2014,53.1,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2014,11.7,"Malta"
"Y15-24","MT0",2014,11.7,"Malta"
"Y15-24","MT00",2014,11.7,"Malta"
"Y15-24","NL",2014,12.7,"Netherlands"
"Y15-24","NL1",2014,14.5,"Noord-Nederland"
"Y15-24","NL11",2014,15.6,"Groningen"
"Y15-24","NL12",2014,13.5,"Friesland (NL)"
"Y15-24","NL13",2014,14.5,"Drenthe"
"Y15-24","NL2",2014,12.3,"Oost-Nederland"
"Y15-24","NL21",2014,12.2,"Overijssel"
"Y15-24","NL22",2014,10.5,"Gelderland"
"Y15-24","NL23",2014,21.2,"Flevoland"
"Y15-24","NL3",2014,12.8,"West-Nederland"
"Y15-24","NL31",2014,11.5,"Utrecht"
"Y15-24","NL32",2014,12,"Noord-Holland"
"Y15-24","NL33",2014,14.3,"Zuid-Holland"
"Y15-24","NL34",2014,9,"Zeeland"
"Y15-24","NL4",2014,12.1,"Zuid-Nederland"
"Y15-24","NL41",2014,11.5,"Noord-Brabant"
"Y15-24","NL42",2014,13.6,"Limburg (NL)"
"Y15-24","NO",2014,7.9,"Norway"
"Y15-24","NO0",2014,7.9,"Norge"
"Y15-24","NO01",2014,7.3,"Oslo og Akershus"
"Y15-24","NO02",2014,6.9,"Hedmark og Oppland"
"Y15-24","NO03",2014,9.7,"Sør-Østlandet"
"Y15-24","NO04",2014,6.5,"Agder og Rogaland"
"Y15-24","NO05",2014,7.4,"Vestlandet"
"Y15-24","NO06",2014,7.7,"Trøndelag"
"Y15-24","NO07",2014,9.7,"Nord-Norge"
"Y15-24","PL",2014,23.9,"Poland"
"Y15-24","PL1",2014,18.5,"Region Centralny"
"Y15-24","PL11",2014,20.1,"Lódzkie"
"Y15-24","PL12",2014,17.7,"Mazowieckie"
"Y15-24","PL2",2014,23.4,"Region Poludniowy"
"Y15-24","PL21",2014,24.8,"Malopolskie"
"Y15-24","PL22",2014,22.2,"Slaskie"
"Y15-24","PL3",2014,33.2,"Region Wschodni"
"Y15-24","PL31",2014,33.2,"Lubelskie"
"Y15-24","PL32",2014,41.1,"Podkarpackie"
"Y15-24","PL33",2014,26.8,"Swietokrzyskie"
"Y15-24","PL34",2014,27,"Podlaskie"
"Y15-24","PL4",2014,22.5,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2014,20.7,"Wielkopolskie"
"Y15-24","PL42",2014,25.1,"Zachodniopomorskie"
"Y15-24","PL43",2014,27.2,"Lubuskie"
"Y15-24","PL5",2014,22.5,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2014,23.5,"Dolnoslaskie"
"Y15-24","PL52",2014,19.9,"Opolskie"
"Y15-24","PL6",2014,24.2,"Region Pólnocny"
"Y15-24","PL61",2014,26.6,"Kujawsko-Pomorskie"
"Y15-24","PL62",2014,25.4,"Warminsko-Mazurskie"
"Y15-24","PL63",2014,21.6,"Pomorskie"
"Y15-24","PT",2014,34.8,"Portugal"
"Y15-24","PT1",2014,34.1,"Continente"
"Y15-24","PT11",2014,35.7,"Norte"
"Y15-24","PT15",2014,30.2,"Algarve"
"Y15-24","PT16",2014,28.2,"Centro (PT)"
"Y15-24","PT17",2014,36.7,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2014,36.2,"Alentejo"
"Y15-24","PT2",2014,41.5,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2014,41.5,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2014,50.5,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2014,50.5,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2014,24,"Romania"
"Y15-24","RO1",2014,22.9,"Macroregiunea unu"
"Y15-24","RO11",2014,13.8,"Nord-Vest"
"Y15-24","RO12",2014,34,"Centru"
"Y15-24","RO2",2014,18.7,"Macroregiunea doi"
"Y15-24","RO21",2014,12.4,"Nord-Est"
"Y15-24","RO22",2014,29.5,"Sud-Est"
"Y15-24","RO3",2014,31.3,"Macroregiunea trei"
"Y15-24","RO31",2014,33.8,"Sud - Muntenia"
"Y15-24","RO32",2014,26.4,"Bucuresti - Ilfov"
"Y15-24","RO4",2014,24.9,"Macroregiunea patru"
"Y15-24","RO41",2014,23.4,"Sud-Vest Oltenia"
"Y15-24","RO42",2014,27.3,"Vest"
"Y15-24","SE",2014,22.9,"Sweden"
"Y15-24","SE1",2014,22.7,"Östra Sverige"
"Y15-24","SE11",2014,21.5,"Stockholm"
"Y15-24","SE12",2014,24.2,"Östra Mellansverige"
"Y15-24","SE2",2014,23.1,"Södra Sverige"
"Y15-24","SE21",2014,19.4,"Småland med öarna"
"Y15-24","SE22",2014,26.1,"Sydsverige"
"Y15-24","SE23",2014,22.7,"Västsverige"
"Y15-24","SE3",2014,22.6,"Norra Sverige"
"Y15-24","SE31",2014,24.5,"Norra Mellansverige"
"Y15-24","SE32",2014,20.3,"Mellersta Norrland"
"Y15-24","SE33",2014,21.3,"Övre Norrland"
"Y15-24","SI",2014,20.2,"Slovenia"
"Y15-24","SI0",2014,20.2,"Slovenija"
"Y15-24","SI03",2014,24,"Vzhodna Slovenija"
"Y15-24","SI04",2014,15.9,"Zahodna Slovenija"
"Y15-24","SK",2014,29.7,"Slovakia"
"Y15-24","SK0",2014,29.7,"Slovensko"
"Y15-24","SK01",2014,14.7,"Bratislavský kraj"
"Y15-24","SK02",2014,25.9,"Západné Slovensko"
"Y15-24","SK03",2014,33.5,"Stredné Slovensko"
"Y15-24","SK04",2014,34.8,"Východné Slovensko"
"Y15-24","TR",2014,17.8,"Turkey"
"Y15-24","TR1",2014,18.9,"Istanbul"
"Y15-24","TR10",2014,18.9,"Istanbul"
"Y15-24","TR2",2014,14.5,"Bati Marmara"
"Y15-24","TR21",2014,13.2,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2014,16.5,"Balikesir, Çanakkale"
"Y15-24","TR3",2014,17,"Ege"
"Y15-24","TR31",2014,22.2,"Izmir"
"Y15-24","TR32",2014,14.4,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2014,10.5,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2014,15.9,"Dogu Marmara"
"Y15-24","TR41",2014,11.3,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2014,20.1,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2014,18.1,"Bati Anadolu"
"Y15-24","TR51",2014,21.6,"Ankara"
"Y15-24","TR52",2014,11.5,"Konya, Karaman"
"Y15-24","TR6",2014,19.5,"Akdeniz"
"Y15-24","TR61",2014,15.6,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2014,17.9,"Adana, Mersin"
"Y15-24","TR63",2014,25.3,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2014,15.9,"Orta Anadolu"
"Y15-24","TR71",2014,13.8,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2014,17,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2014,13.6,"Bati Karadeniz"
"Y15-24","TR81",2014,15.2,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2014,16.6,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2014,12.1,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2014,18.4,"Dogu Karadeniz"
"Y15-24","TR90",2014,18.4,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2014,9.2,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2014,13.5,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2014,5.9,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2014,18.7,"Ortadogu Anadolu"
"Y15-24","TRB1",2014,15,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2014,20.7,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2014,21.9,"Güneydogu Anadolu"
"Y15-24","TRC1",2014,16.1,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2014,19.5,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2014,33.1,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2014,17,"United Kingdom"
"Y15-24","UKC",2014,23,"North East (UK)"
"Y15-24","UKC1",2014,24.8,"Tees Valley and Durham"
"Y15-24","UKC2",2014,21.5,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2014,16.5,"North West (UK)"
"Y15-24","UKD1",2014,11,"Cumbria"
"Y15-24","UKD3",2014,18.5,"Greater Manchester"
"Y15-24","UKD4",2014,15,"Lancashire"
"Y15-24","UKD6",2014,9.1,"Cheshire"
"Y15-24","UKD7",2014,20.2,"Merseyside"
"Y15-24","UKE",2014,17.8,"Yorkshire and The Humber"
"Y15-24","UKE1",2014,17.5,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2014,12.5,"North Yorkshire"
"Y15-24","UKE3",2014,20.3,"South Yorkshire"
"Y15-24","UKE4",2014,17.7,"West Yorkshire"
"Y15-24","UKF",2014,13.2,"East Midlands (UK)"
"Y15-24","UKF1",2014,16,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2014,11.8,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2014,8.6,"Lincolnshire"
"Y15-24","UKG",2014,20,"West Midlands (UK)"
"Y15-24","UKG1",2014,13.1,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2014,13.4,"Shropshire and Staffordshire"
"Y15-24","UKG3",2014,26.8,"West Midlands"
"Y15-24","UKH",2014,15.2,"East of England"
"Y15-24","UKH1",2014,14.5,"East Anglia"
"Y15-24","UKH2",2014,15.2,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2014,16.3,"Essex"
"Y15-24","UKI",2014,19.4,"London"
"Y15-24","UKI3",2014,11.6,"Inner London - West"
"Y15-24","UKI4",2014,21.6,"Inner London - East"
"Y15-24","UKI5",2014,21.9,"Outer London - East and North East"
"Y15-24","UKI6",2014,18.3,"Outer London - South"
"Y15-24","UKI7",2014,19.8,"Outer London - West and North West"
"Y15-24","UKJ",2014,14.9,"South East (UK)"
"Y15-24","UKJ1",2014,13.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2014,16.6,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2014,13.2,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2014,16.3,"Kent"
"Y15-24","UKK",2014,14.2,"South West (UK)"
"Y15-24","UKK1",2014,12.6,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2014,16.3,"Dorset and Somerset"
"Y15-24","UKK3",2014,11.2,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2014,17,"Devon"
"Y15-24","UKL",2014,18.6,"Wales"
"Y15-24","UKL1",2014,18.8,"West Wales and The Valleys"
"Y15-24","UKL2",2014,18.2,"East Wales"
"Y15-24","UKM",2014,16.7,"Scotland"
"Y15-24","UKM2",2014,17.5,"Eastern Scotland"
"Y15-24","UKM3",2014,19.3,"South Western Scotland"
"Y15-24","UKM5",2014,NA,"North Eastern Scotland"
"Y15-24","UKM6",2014,14.5,"Highlands and Islands"
"Y15-24","UKN",2014,19.7,"Northern Ireland (UK)"
"Y15-24","UKN0",2014,19.7,"Northern Ireland (UK)"
"Y20-64","AT",2014,5.5,"Austria"
"Y20-64","AT1",2014,7.2,"Ostösterreich"
"Y20-64","AT11",2014,4.7,"Burgenland (AT)"
"Y20-64","AT12",2014,4.7,"Niederösterreich"
"Y20-64","AT13",2014,9.9,"Wien"
"Y20-64","AT2",2014,5.2,"Südösterreich"
"Y20-64","AT21",2014,5.8,"Kärnten"
"Y20-64","AT22",2014,5,"Steiermark"
"Y20-64","AT3",2014,3.6,"Westösterreich"
"Y20-64","AT31",2014,4,"Oberösterreich"
"Y20-64","AT32",2014,3.5,"Salzburg"
"Y20-64","AT33",2014,3.1,"Tirol"
"Y20-64","AT34",2014,3.1,"Vorarlberg"
"Y20-64","BE",2014,8.4,"Belgium"
"Y20-64","BE1",2014,18.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2014,18.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2014,4.9,"Vlaams Gewest"
"Y20-64","BE21",2014,5.9,"Prov. Antwerpen"
"Y20-64","BE22",2014,5.4,"Prov. Limburg (BE)"
"Y20-64","BE23",2014,4.1,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2014,4.8,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2014,4,"Prov. West-Vlaanderen"
"Y20-64","BE3",2014,11.7,"Région wallonne"
"Y20-64","BE31",2014,8.6,"Prov. Brabant Wallon"
"Y20-64","BE32",2014,14.2,"Prov. Hainaut"
"Y20-64","BE33",2014,12.3,"Prov. Liège"
"Y20-64","BE34",2014,8.4,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2014,8.8,"Prov. Namur"
"Y20-64","BG",2014,11.3,"Bulgaria"
"Y20-64","BG3",2014,12.8,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2014,14.1,"Severozapaden"
"Y20-64","BG32",2014,13.1,"Severen tsentralen"
"Y20-64","BG33",2014,12.6,"Severoiztochen"
"Y20-64","BG34",2014,11.8,"Yugoiztochen"
"Y20-64","BG4",2014,10,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2014,8.9,"Yugozapaden"
"Y20-64","BG42",2014,11.9,"Yuzhen tsentralen"
"Y20-64","CH",2014,4.5,"Switzerland"
"Y20-64","CH0",2014,4.5,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2014,6.4,"Région lémanique"
"Y20-64","CH02",2014,4.2,"Espace Mittelland"
"Y20-64","CH03",2014,4.3,"Nordwestschweiz"
"Y20-64","CH04",2014,4.2,"Zürich"
"Y20-64","CH05",2014,3.2,"Ostschweiz"
"Y20-64","CH06",2014,3.5,"Zentralschweiz"
"Y20-64","CH07",2014,6.7,"Ticino"
"Y20-64","CY",2014,16,"Cyprus"
"Y20-64","CY0",2014,16,"Kypros"
"Y20-64","CY00",2014,16,"Kypros"
"Y20-64","CZ",2014,6,"Czech Republic"
"Y20-64","CZ0",2014,6,"Ceská republika"
"Y20-64","CZ01",2014,2.4,"Praha"
"Y20-64","CZ02",2014,5.1,"Strední Cechy"
"Y20-64","CZ03",2014,5.4,"Jihozápad"
"Y20-64","CZ04",2014,8.5,"Severozápad"
"Y20-64","CZ05",2014,6.2,"Severovýchod"
"Y20-64","CZ06",2014,5.8,"Jihovýchod"
"Y20-64","CZ07",2014,6.7,"Strední Morava"
"Y20-64","CZ08",2014,8.5,"Moravskoslezsko"
"Y20-64","DE",2014,5,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2014,3.1,"Baden-Württemberg"
"Y20-64","DE11",2014,3.1,"Stuttgart"
"Y20-64","DE12",2014,3.5,"Karlsruhe"
"Y20-64","DE13",2014,3,"Freiburg"
"Y20-64","DE14",2014,2.5,"Tübingen"
"Y20-64","DE2",2014,2.8,"Bayern"
"Y20-64","DE21",2014,2.5,"Oberbayern"
"Y20-64","DE22",2014,2.8,"Niederbayern"
"Y20-64","DE23",2014,2.8,"Oberpfalz"
"Y20-64","DE24",2014,3.9,"Oberfranken"
"Y20-64","DE25",2014,3.1,"Mittelfranken"
"Y20-64","DE26",2014,2.9,"Unterfranken"
"Y20-64","DE27",2014,2.9,"Schwaben"
"Y20-64","DE3",2014,9.8,"Berlin"
"Y20-64","DE30",2014,9.8,"Berlin"
"Y20-64","DE4",2014,6.7,"Brandenburg"
"Y20-64","DE40",2014,6.7,"Brandenburg"
"Y20-64","DE5",2014,6.5,"Bremen"
"Y20-64","DE50",2014,6.5,"Bremen"
"Y20-64","DE6",2014,4.9,"Hamburg"
"Y20-64","DE60",2014,4.9,"Hamburg"
"Y20-64","DE7",2014,4.3,"Hessen"
"Y20-64","DE71",2014,4.3,"Darmstadt"
"Y20-64","DE72",2014,4.1,"Gießen"
"Y20-64","DE73",2014,4.3,"Kassel"
"Y20-64","DE8",2014,9.7,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2014,9.7,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2014,4.6,"Niedersachsen"
"Y20-64","DE91",2014,5.4,"Braunschweig"
"Y20-64","DE92",2014,5.2,"Hannover"
"Y20-64","DE93",2014,4,"Lüneburg"
"Y20-64","DE94",2014,4.1,"Weser-Ems"
"Y20-64","DEA",2014,5.6,"Nordrhein-Westfalen"
"Y20-64","DEA1",2014,6.3,"Düsseldorf"
"Y20-64","DEA2",2014,5.2,"Köln"
"Y20-64","DEA3",2014,4.9,"Münster"
"Y20-64","DEA4",2014,5,"Detmold"
"Y20-64","DEA5",2014,5.7,"Arnsberg"
"Y20-64","DEB",2014,3.8,"Rheinland-Pfalz"
"Y20-64","DEB1",2014,4,"Koblenz"
"Y20-64","DEB2",2014,2.7,"Trier"
"Y20-64","DEB3",2014,3.9,"Rheinhessen-Pfalz"
"Y20-64","DEC",2014,5.9,"Saarland"
"Y20-64","DEC0",2014,5.9,"Saarland"
"Y20-64","DED",2014,7.3,"Sachsen"
"Y20-64","DED2",2014,7.3,"Dresden"
"Y20-64","DED4",2014,6.5,"Chemnitz"
"Y20-64","DED5",2014,8.3,"Leipzig"
"Y20-64","DEE",2014,8.8,"Sachsen-Anhalt"
"Y20-64","DEE0",2014,8.8,"Sachsen-Anhalt"
"Y20-64","DEF",2014,4.5,"Schleswig-Holstein"
"Y20-64","DEF0",2014,4.5,"Schleswig-Holstein"
"Y20-64","DEG",2014,6,"Thüringen"
"Y20-64","DEG0",2014,6,"Thüringen"
"Y20-64","DK",2014,6.2,"Denmark"
"Y20-64","DK0",2014,6.2,"Danmark"
"Y20-64","DK01",2014,6.7,"Hovedstaden"
"Y20-64","DK02",2014,5.8,"Sjælland"
"Y20-64","DK03",2014,6.3,"Syddanmark"
"Y20-64","DK04",2014,5.8,"Midtjylland"
"Y20-64","DK05",2014,6.1,"Nordjylland"
"Y20-64","EA17",2014,11.5,"Euro area (17 countries)"
"Y20-64","EA18",2014,11.5,"Euro area (18 countries)"
"Y20-64","EA19",2014,11.5,"Euro area (19 countries)"
"Y20-64","EE",2014,7.3,"Estonia"
"Y20-64","EE0",2014,7.3,"Eesti"
"Y20-64","EE00",2014,7.3,"Eesti"
"Y20-64","EL",2014,26.4,"Greece"
"Y20-64","EL3",2014,27.2,"Attiki"
"Y20-64","EL30",2014,27.2,"Attiki"
"Y20-64","EL4",2014,22.5,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2014,22.3,"Voreio Aigaio"
"Y20-64","EL42",2014,20.4,"Notio Aigaio"
"Y20-64","EL43",2014,23.8,"Kriti"
"Y20-64","EL5",2014,27.4,"Voreia Ellada"
"Y20-64","EL51",2014,23.9,"Anatoliki Makedonia, Thraki"
"Y20-64","EL52",2014,28.6,"Kentriki Makedonia"
"Y20-64","EL53",2014,27.4,"Dytiki Makedonia"
"Y20-64","EL54",2014,27,"Ipeiros"
"Y20-64","EL6",2014,25.8,"Kentriki Ellada"
"Y20-64","EL61",2014,25.9,"Thessalia"
"Y20-64","EL62",2014,21.2,"Ionia Nisia"
"Y20-64","EL63",2014,28.5,"Dytiki Ellada"
"Y20-64","EL64",2014,26.8,"Sterea Ellada"
"Y20-64","EL65",2014,23.4,"Peloponnisos"
"Y20-64","ES",2014,24.1,"Spain"
"Y20-64","ES1",2014,21.1,"Noroeste (ES)"
"Y20-64","ES11",2014,21.5,"Galicia"
"Y20-64","ES12",2014,21,"Principado de Asturias"
"Y20-64","ES13",2014,19.4,"Cantabria"
"Y20-64","ES2",2014,17.2,"Noreste (ES)"
"Y20-64","ES21",2014,16.2,"País Vasco"
"Y20-64","ES22",2014,15.1,"Comunidad Foral de Navarra"
"Y20-64","ES23",2014,17.7,"La Rioja"
"Y20-64","ES24",2014,19.8,"Aragón"
"Y20-64","ES3",2014,18.3,"Comunidad de Madrid"
"Y20-64","ES30",2014,18.3,"Comunidad de Madrid"
"Y20-64","ES4",2014,25.1,"Centro (ES)"
"Y20-64","ES41",2014,20.5,"Castilla y León"
"Y20-64","ES42",2014,28.4,"Castilla-la Mancha"
"Y20-64","ES43",2014,29.3,"Extremadura"
"Y20-64","ES5",2014,21.8,"Este (ES)"
"Y20-64","ES51",2014,19.9,"Cataluña"
"Y20-64","ES52",2014,25.4,"Comunidad Valenciana"
"Y20-64","ES53",2014,19.5,"Illes Balears"
"Y20-64","ES6",2014,33.1,"Sur (ES)"
"Y20-64","ES61",2014,34.4,"Andalucía"
"Y20-64","ES62",2014,26.2,"Región de Murcia"
"Y20-64","ES63",2014,31.1,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2014,28,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2014,32.2,"Canarias (ES)"
"Y20-64","ES70",2014,32.2,"Canarias (ES)"
"Y20-64","EU15",2014,10.3,"European Union (15 countries)"
"Y20-64","EU27",2014,10,"European Union (27 countries)"
"Y20-64","EU28",2014,10,"European Union (28 countries)"
"Y20-64","FI",2014,8,"Finland"
"Y20-64","FI1",2014,8.1,"Manner-Suomi"
"Y20-64","FI19",2014,8.2,"Länsi-Suomi"
"Y20-64","FI1B",2014,6.7,"Helsinki-Uusimaa"
"Y20-64","FI1C",2014,8.7,"Etelä-Suomi"
"Y20-64","FI1D",2014,9.3,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2014,NA,"Åland"
"Y20-64","FI20",2014,NA,"Åland"
"Y20-64","FR",2014,9.9,"France"
"Y20-64","FR1",2014,9.5,"Île de France"
"Y20-64","FR10",2014,9.5,"Île de France"
"Y20-64","FR2",2014,10.2,"Bassin Parisien"
"Y20-64","FR21",2014,11.1,"Champagne-Ardenne"
"Y20-64","FR22",2014,11,"Picardie"
"Y20-64","FR23",2014,11.4,"Haute-Normandie"
"Y20-64","FR24",2014,9.2,"Centre (FR)"
"Y20-64","FR25",2014,7.9,"Basse-Normandie"
"Y20-64","FR26",2014,10.4,"Bourgogne"
"Y20-64","FR3",2014,13.2,"Nord - Pas-de-Calais"
"Y20-64","FR30",2014,13.2,"Nord - Pas-de-Calais"
"Y20-64","FR4",2014,10.3,"Est (FR)"
"Y20-64","FR41",2014,11.4,"Lorraine"
"Y20-64","FR42",2014,9.4,"Alsace"
"Y20-64","FR43",2014,9.5,"Franche-Comté"
"Y20-64","FR5",2014,8.2,"Ouest (FR)"
"Y20-64","FR51",2014,8.2,"Pays de la Loire"
"Y20-64","FR52",2014,7.1,"Bretagne"
"Y20-64","FR53",2014,10.4,"Poitou-Charentes"
"Y20-64","FR6",2014,8.7,"Sud-Ouest (FR)"
"Y20-64","FR61",2014,8.6,"Aquitaine"
"Y20-64","FR62",2014,8.7,"Midi-Pyrénées"
"Y20-64","FR63",2014,8.9,"Limousin"
"Y20-64","FR7",2014,8.2,"Centre-Est (FR)"
"Y20-64","FR71",2014,8.4,"Rhône-Alpes"
"Y20-64","FR72",2014,7,"Auvergne"
"Y20-64","FR8",2014,10.4,"Méditerranée"
"Y20-64","FR81",2014,11.8,"Languedoc-Roussillon"
"Y20-64","FR82",2014,9.7,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2014,9.3,"Corse"
"Y20-64","FRA",2014,23.1,"Départements d'outre-mer"
"Y20-64","FRA1",2014,23.6,"Guadeloupe"
"Y20-64","FRA2",2014,19,"Martinique"
"Y20-64","FRA3",2014,21.8,"Guyane"
"Y20-64","FRA4",2014,25.7,"La Réunion"
"Y20-64","FRA5",2014,19,"Mayotte"
"Y20-64","HR",2014,16.5,"Croatia"
"Y20-64","HR0",2014,16.5,"Hrvatska"
"Y20-64","HR03",2014,16.3,"Jadranska Hrvatska"
"Y20-64","HR04",2014,16.7,"Kontinentalna Hrvatska"
"Y20-64","HU",2014,7.6,"Hungary"
"Y20-64","HU1",2014,6.1,"Közép-Magyarország"
"Y20-64","HU10",2014,6.1,"Közép-Magyarország"
"Y20-64","HU2",2014,5.7,"Dunántúl"
"Y20-64","HU21",2014,5.4,"Közép-Dunántúl"
"Y20-64","HU22",2014,4.4,"Nyugat-Dunántúl"
"Y20-64","HU23",2014,7.6,"Dél-Dunántúl"
"Y20-64","HU3",2014,10.3,"Alföld és Észak"
"Y20-64","HU31",2014,10.2,"Észak-Magyarország"
"Y20-64","HU32",2014,11.5,"Észak-Alföld"
"Y20-64","HU33",2014,8.8,"Dél-Alföld"
"Y20-64","IE",2014,11.1,"Ireland"
"Y20-64","IE0",2014,11.1,"Éire/Ireland"
"Y20-64","IE01",2014,12.3,"Border, Midland and Western"
"Y20-64","IE02",2014,10.7,"Southern and Eastern"
"Y20-64","IS",2014,4.4,"Iceland"
"Y20-64","IS0",2014,4.4,"Ísland"
"Y20-64","IS00",2014,4.4,"Ísland"
"Y20-64","IT",2014,12.5,"Italy"
"Y20-64","ITC",2014,9.1,"Nord-Ovest"
"Y20-64","ITC1",2014,11.1,"Piemonte"
"Y20-64","ITC2",2014,8.7,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2014,10.7,"Liguria"
"Y20-64","ITC4",2014,7.9,"Lombardia"
"Y20-64","ITF",2014,20,"Sud"
"Y20-64","ITF1",2014,12.6,"Abruzzo"
"Y20-64","ITF2",2014,15,"Molise"
"Y20-64","ITF3",2014,21.3,"Campania"
"Y20-64","ITF4",2014,20.9,"Puglia"
"Y20-64","ITF5",2014,14.6,"Basilicata"
"Y20-64","ITF6",2014,23.1,"Calabria"
"Y20-64","ITG",2014,20.9,"Isole"
"Y20-64","ITG1",2014,21.8,"Sicilia"
"Y20-64","ITG2",2014,18.5,"Sardegna"
"Y20-64","ITH",2014,7.5,"Nord-Est"
"Y20-64","ITH1",2014,4.2,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2014,6.8,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2014,7.2,"Veneto"
"Y20-64","ITH4",2014,8,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2014,8.2,"Emilia-Romagna"
"Y20-64","ITI",2014,11.3,"Centro (IT)"
"Y20-64","ITI1",2014,10,"Toscana"
"Y20-64","ITI2",2014,11.2,"Umbria"
"Y20-64","ITI3",2014,9.9,"Marche"
"Y20-64","ITI4",2014,12.4,"Lazio"
"Y20-64","LT",2014,10.8,"Lithuania"
"Y20-64","LT0",2014,10.8,"Lietuva"
"Y20-64","LT00",2014,10.8,"Lietuva"
"Y20-64","LU",2014,5.6,"Luxembourg"
"Y20-64","LU0",2014,5.6,"Luxembourg"
"Y20-64","LU00",2014,5.6,"Luxembourg"
"Y20-64","LV",2014,10.9,"Latvia"
"Y20-64","LV0",2014,10.9,"Latvija"
"Y20-64","LV00",2014,10.9,"Latvija"
"Y20-64","MK",2014,27.5,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2014,27.5,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2014,27.5,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2014,5.3,"Malta"
"Y20-64","MT0",2014,5.3,"Malta"
"Y20-64","MT00",2014,5.3,"Malta"
"Y20-64","NL",2014,6.9,"Netherlands"
"Y20-64","NL1",2014,7.4,"Noord-Nederland"
"Y20-64","NL11",2014,7.9,"Groningen"
"Y20-64","NL12",2014,7.4,"Friesland (NL)"
"Y20-64","NL13",2014,6.6,"Drenthe"
"Y20-64","NL2",2014,7,"Oost-Nederland"
"Y20-64","NL21",2014,6.6,"Overijssel"
"Y20-64","NL22",2014,6.6,"Gelderland"
"Y20-64","NL23",2014,10,"Flevoland"
"Y20-64","NL3",2014,6.9,"West-Nederland"
"Y20-64","NL31",2014,5.9,"Utrecht"
"Y20-64","NL32",2014,6.3,"Noord-Holland"
"Y20-64","NL33",2014,7.9,"Zuid-Holland"
"Y20-64","NL34",2014,4.5,"Zeeland"
"Y20-64","NL4",2014,6.5,"Zuid-Nederland"
"Y20-64","NL41",2014,6.5,"Noord-Brabant"
"Y20-64","NL42",2014,6.8,"Limburg (NL)"
"Y20-64","NO",2014,3.3,"Norway"
"Y20-64","NO0",2014,3.3,"Norge"
"Y20-64","NO01",2014,3.7,"Oslo og Akershus"
"Y20-64","NO02",2014,2.6,"Hedmark og Oppland"
"Y20-64","NO03",2014,3.8,"Sør-Østlandet"
"Y20-64","NO04",2014,2.8,"Agder og Rogaland"
"Y20-64","NO05",2014,2.7,"Vestlandet"
"Y20-64","NO06",2014,3.6,"Trøndelag"
"Y20-64","NO07",2014,2.9,"Nord-Norge"
"Y20-64","PL",2014,8.9,"Poland"
"Y20-64","PL1",2014,7.7,"Region Centralny"
"Y20-64","PL11",2014,8.9,"Lódzkie"
"Y20-64","PL12",2014,7.1,"Mazowieckie"
"Y20-64","PL2",2014,8.7,"Region Poludniowy"
"Y20-64","PL21",2014,9,"Malopolskie"
"Y20-64","PL22",2014,8.5,"Slaskie"
"Y20-64","PL3",2014,11.3,"Region Wschodni"
"Y20-64","PL31",2014,9.9,"Lubelskie"
"Y20-64","PL32",2014,14,"Podkarpackie"
"Y20-64","PL33",2014,11.5,"Swietokrzyskie"
"Y20-64","PL34",2014,9.1,"Podlaskie"
"Y20-64","PL4",2014,7.8,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2014,7.5,"Wielkopolskie"
"Y20-64","PL42",2014,8.3,"Zachodniopomorskie"
"Y20-64","PL43",2014,8.2,"Lubuskie"
"Y20-64","PL5",2014,8.8,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2014,9.1,"Dolnoslaskie"
"Y20-64","PL52",2014,7.7,"Opolskie"
"Y20-64","PL6",2014,9.5,"Region Pólnocny"
"Y20-64","PL61",2014,10.5,"Kujawsko-Pomorskie"
"Y20-64","PL62",2014,9.6,"Warminsko-Mazurskie"
"Y20-64","PL63",2014,8.5,"Pomorskie"
"Y20-64","PT",2014,14.1,"Portugal"
"Y20-64","PT1",2014,14,"Continente"
"Y20-64","PT11",2014,15,"Norte"
"Y20-64","PT15",2014,14.5,"Algarve"
"Y20-64","PT16",2014,11.1,"Centro (PT)"
"Y20-64","PT17",2014,14.8,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2014,14.5,"Alentejo"
"Y20-64","PT2",2014,15.9,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2014,15.9,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2014,15.4,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2014,15.4,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2014,6.7,"Romania"
"Y20-64","RO1",2014,6,"Macroregiunea unu"
"Y20-64","RO11",2014,3.8,"Nord-Vest"
"Y20-64","RO12",2014,8.7,"Centru"
"Y20-64","RO2",2014,6.6,"Macroregiunea doi"
"Y20-64","RO21",2014,4.3,"Nord-Est"
"Y20-64","RO22",2014,10,"Sud-Est"
"Y20-64","RO3",2014,8,"Macroregiunea trei"
"Y20-64","RO31",2014,8.8,"Sud - Muntenia"
"Y20-64","RO32",2014,6.9,"Bucuresti - Ilfov"
"Y20-64","RO4",2014,5.8,"Macroregiunea patru"
"Y20-64","RO41",2014,6.8,"Sud-Vest Oltenia"
"Y20-64","RO42",2014,4.6,"Vest"
"Y20-64","SE",2014,7.1,"Sweden"
"Y20-64","SE1",2014,6.7,"Östra Sverige"
"Y20-64","SE11",2014,6.2,"Stockholm"
"Y20-64","SE12",2014,7.4,"Östra Mellansverige"
"Y20-64","SE2",2014,7.4,"Södra Sverige"
"Y20-64","SE21",2014,6,"Småland med öarna"
"Y20-64","SE22",2014,9.1,"Sydsverige"
"Y20-64","SE23",2014,6.7,"Västsverige"
"Y20-64","SE3",2014,7.2,"Norra Sverige"
"Y20-64","SE31",2014,7.9,"Norra Mellansverige"
"Y20-64","SE32",2014,6.7,"Mellersta Norrland"
"Y20-64","SE33",2014,6.5,"Övre Norrland"
"Y20-64","SI",2014,9.8,"Slovenia"
"Y20-64","SI0",2014,9.8,"Slovenija"
"Y20-64","SI03",2014,11.2,"Vzhodna Slovenija"
"Y20-64","SI04",2014,8.2,"Zahodna Slovenija"
"Y20-64","SK",2014,12.9,"Slovakia"
"Y20-64","SK0",2014,12.9,"Slovensko"
"Y20-64","SK01",2014,5.9,"Bratislavský kraj"
"Y20-64","SK02",2014,10.7,"Západné Slovensko"
"Y20-64","SK03",2014,15.7,"Stredné Slovensko"
"Y20-64","SK04",2014,16.2,"Východné Slovensko"
"Y20-64","TR",2014,9.7,"Turkey"
"Y20-64","TR1",2014,11.4,"Istanbul"
"Y20-64","TR10",2014,11.4,"Istanbul"
"Y20-64","TR2",2014,6.7,"Bati Marmara"
"Y20-64","TR21",2014,7.7,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2014,5.6,"Balikesir, Çanakkale"
"Y20-64","TR3",2014,8.9,"Ege"
"Y20-64","TR31",2014,13.3,"Izmir"
"Y20-64","TR32",2014,7.4,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2014,3.9,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2014,7.8,"Dogu Marmara"
"Y20-64","TR41",2014,6,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2014,9.6,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2014,9.5,"Bati Anadolu"
"Y20-64","TR51",2014,11.1,"Ankara"
"Y20-64","TR52",2014,5.5,"Konya, Karaman"
"Y20-64","TR6",2014,11,"Akdeniz"
"Y20-64","TR61",2014,8.3,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2014,10.8,"Adana, Mersin"
"Y20-64","TR63",2014,14.8,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2014,8.7,"Orta Anadolu"
"Y20-64","TR71",2014,7.7,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2014,9.3,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2014,6.3,"Bati Karadeniz"
"Y20-64","TR81",2014,6.1,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2014,6.6,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2014,6.3,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2014,6.4,"Dogu Karadeniz"
"Y20-64","TR90",2014,6.4,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2014,5.3,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2014,7.4,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2014,3.3,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2014,10.3,"Ortadogu Anadolu"
"Y20-64","TRB1",2014,7.4,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2014,13,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2014,15.3,"Güneydogu Anadolu"
"Y20-64","TRC1",2014,7.5,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2014,17.9,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2014,23,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2014,5.4,"United Kingdom"
"Y20-64","UKC",2014,7.9,"North East (UK)"
"Y20-64","UKC1",2014,8.5,"Tees Valley and Durham"
"Y20-64","UKC2",2014,7.5,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2014,5.8,"North West (UK)"
"Y20-64","UKD1",2014,4.3,"Cumbria"
"Y20-64","UKD3",2014,6.9,"Greater Manchester"
"Y20-64","UKD4",2014,5.8,"Lancashire"
"Y20-64","UKD6",2014,2.9,"Cheshire"
"Y20-64","UKD7",2014,6.3,"Merseyside"
"Y20-64","UKE",2014,6.3,"Yorkshire and The Humber"
"Y20-64","UKE1",2014,7.4,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2014,3.8,"North Yorkshire"
"Y20-64","UKE3",2014,7.5,"South Yorkshire"
"Y20-64","UKE4",2014,6,"West Yorkshire"
"Y20-64","UKF",2014,5,"East Midlands (UK)"
"Y20-64","UKF1",2014,5.5,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2014,4.8,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2014,4.4,"Lincolnshire"
"Y20-64","UKG",2014,6.3,"West Midlands (UK)"
"Y20-64","UKG1",2014,3.6,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2014,4.8,"Shropshire and Staffordshire"
"Y20-64","UKG3",2014,8.5,"West Midlands"
"Y20-64","UKH",2014,4.5,"East of England"
"Y20-64","UKH1",2014,4.2,"East Anglia"
"Y20-64","UKH2",2014,3.8,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2014,5.6,"Essex"
"Y20-64","UKI",2014,6.1,"London"
"Y20-64","UKI3",2014,5.6,"Inner London - West"
"Y20-64","UKI4",2014,7.1,"Inner London - East"
"Y20-64","UKI5",2014,6.7,"Outer London - East and North East"
"Y20-64","UKI6",2014,4.8,"Outer London - South"
"Y20-64","UKI7",2014,5.3,"Outer London - West and North West"
"Y20-64","UKJ",2014,3.9,"South East (UK)"
"Y20-64","UKJ1",2014,3.7,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2014,3.8,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2014,3.6,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2014,4.9,"Kent"
"Y20-64","UKK",2014,4,"South West (UK)"
"Y20-64","UKK1",2014,4.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2014,3.7,"Dorset and Somerset"
"Y20-64","UKK3",2014,3.1,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2014,4,"Devon"
"Y20-64","UKL",2014,5.9,"Wales"
"Y20-64","UKL1",2014,6.1,"West Wales and The Valleys"
"Y20-64","UKL2",2014,5.5,"East Wales"
"Y20-64","UKM",2014,5.1,"Scotland"
"Y20-64","UKM2",2014,4.7,"Eastern Scotland"
"Y20-64","UKM3",2014,6.1,"South Western Scotland"
"Y20-64","UKM5",2014,3.7,"North Eastern Scotland"
"Y20-64","UKM6",2014,4.5,"Highlands and Islands"
"Y20-64","UKN",2014,5.8,"Northern Ireland (UK)"
"Y20-64","UKN0",2014,5.8,"Northern Ireland (UK)"
"Y_GE15","AT",2014,5.6,"Austria"
"Y_GE15","AT1",2014,7.5,"Ostösterreich"
"Y_GE15","AT11",2014,4.8,"Burgenland (AT)"
"Y_GE15","AT12",2014,5.1,"Niederösterreich"
"Y_GE15","AT13",2014,10.2,"Wien"
"Y_GE15","AT2",2014,5.2,"Südösterreich"
"Y_GE15","AT21",2014,6,"Kärnten"
"Y_GE15","AT22",2014,4.9,"Steiermark"
"Y_GE15","AT3",2014,3.7,"Westösterreich"
"Y_GE15","AT31",2014,4,"Oberösterreich"
"Y_GE15","AT32",2014,3.5,"Salzburg"
"Y_GE15","AT33",2014,3.2,"Tirol"
"Y_GE15","AT34",2014,3.4,"Vorarlberg"
"Y_GE15","BE",2014,8.5,"Belgium"
"Y_GE15","BE1",2014,18.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2014,18.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2014,5.1,"Vlaams Gewest"
"Y_GE15","BE21",2014,6.1,"Prov. Antwerpen"
"Y_GE15","BE22",2014,5.6,"Prov. Limburg (BE)"
"Y_GE15","BE23",2014,4.3,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2014,5,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2014,4.2,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2014,11.8,"Région wallonne"
"Y_GE15","BE31",2014,8.8,"Prov. Brabant Wallon"
"Y_GE15","BE32",2014,14.4,"Prov. Hainaut"
"Y_GE15","BE33",2014,12.3,"Prov. Liège"
"Y_GE15","BE34",2014,8.5,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2014,8.9,"Prov. Namur"
"Y_GE15","BG",2014,11.4,"Bulgaria"
"Y_GE15","BG3",2014,12.9,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2014,14.2,"Severozapaden"
"Y_GE15","BG32",2014,13.2,"Severen tsentralen"
"Y_GE15","BG33",2014,12.6,"Severoiztochen"
"Y_GE15","BG34",2014,11.9,"Yugoiztochen"
"Y_GE15","BG4",2014,10.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2014,8.9,"Yugozapaden"
"Y_GE15","BG42",2014,12,"Yuzhen tsentralen"
"Y_GE15","CH",2014,4.5,"Switzerland"
"Y_GE15","CH0",2014,4.5,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2014,6.7,"Région lémanique"
"Y_GE15","CH02",2014,4.3,"Espace Mittelland"
"Y_GE15","CH03",2014,4.3,"Nordwestschweiz"
"Y_GE15","CH04",2014,4.1,"Zürich"
"Y_GE15","CH05",2014,3.2,"Ostschweiz"
"Y_GE15","CH06",2014,3.5,"Zentralschweiz"
"Y_GE15","CH07",2014,6.7,"Ticino"
"Y_GE15","CY",2014,16.1,"Cyprus"
"Y_GE15","CY0",2014,16.1,"Kypros"
"Y_GE15","CY00",2014,16.1,"Kypros"
"Y_GE15","CZ",2014,6.1,"Czech Republic"
"Y_GE15","CZ0",2014,6.1,"Ceská republika"
"Y_GE15","CZ01",2014,2.5,"Praha"
"Y_GE15","CZ02",2014,5.1,"Strední Cechy"
"Y_GE15","CZ03",2014,5.5,"Jihozápad"
"Y_GE15","CZ04",2014,8.7,"Severozápad"
"Y_GE15","CZ05",2014,6.3,"Severovýchod"
"Y_GE15","CZ06",2014,5.9,"Jihovýchod"
"Y_GE15","CZ07",2014,6.9,"Strední Morava"
"Y_GE15","CZ08",2014,8.6,"Moravskoslezsko"
"Y_GE15","DE",2014,5,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2014,3.1,"Baden-Württemberg"
"Y_GE15","DE11",2014,3.1,"Stuttgart"
"Y_GE15","DE12",2014,3.5,"Karlsruhe"
"Y_GE15","DE13",2014,3,"Freiburg"
"Y_GE15","DE14",2014,2.6,"Tübingen"
"Y_GE15","DE2",2014,2.9,"Bayern"
"Y_GE15","DE21",2014,2.5,"Oberbayern"
"Y_GE15","DE22",2014,2.8,"Niederbayern"
"Y_GE15","DE23",2014,2.7,"Oberpfalz"
"Y_GE15","DE24",2014,4,"Oberfranken"
"Y_GE15","DE25",2014,3.1,"Mittelfranken"
"Y_GE15","DE26",2014,2.9,"Unterfranken"
"Y_GE15","DE27",2014,3,"Schwaben"
"Y_GE15","DE3",2014,9.8,"Berlin"
"Y_GE15","DE30",2014,9.8,"Berlin"
"Y_GE15","DE4",2014,6.7,"Brandenburg"
"Y_GE15","DE40",2014,6.7,"Brandenburg"
"Y_GE15","DE5",2014,6.6,"Bremen"
"Y_GE15","DE50",2014,6.6,"Bremen"
"Y_GE15","DE6",2014,5,"Hamburg"
"Y_GE15","DE60",2014,5,"Hamburg"
"Y_GE15","DE7",2014,4.4,"Hessen"
"Y_GE15","DE71",2014,4.5,"Darmstadt"
"Y_GE15","DE72",2014,4.5,"Gießen"
"Y_GE15","DE73",2014,4.4,"Kassel"
"Y_GE15","DE8",2014,9.6,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2014,9.6,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2014,4.6,"Niedersachsen"
"Y_GE15","DE91",2014,5.5,"Braunschweig"
"Y_GE15","DE92",2014,5.2,"Hannover"
"Y_GE15","DE93",2014,4,"Lüneburg"
"Y_GE15","DE94",2014,4.1,"Weser-Ems"
"Y_GE15","DEA",2014,5.6,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2014,6.3,"Düsseldorf"
"Y_GE15","DEA2",2014,5.3,"Köln"
"Y_GE15","DEA3",2014,4.9,"Münster"
"Y_GE15","DEA4",2014,5,"Detmold"
"Y_GE15","DEA5",2014,5.7,"Arnsberg"
"Y_GE15","DEB",2014,3.9,"Rheinland-Pfalz"
"Y_GE15","DEB1",2014,4,"Koblenz"
"Y_GE15","DEB2",2014,3,"Trier"
"Y_GE15","DEB3",2014,3.9,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2014,5.8,"Saarland"
"Y_GE15","DEC0",2014,5.8,"Saarland"
"Y_GE15","DED",2014,7.2,"Sachsen"
"Y_GE15","DED2",2014,7.4,"Dresden"
"Y_GE15","DED4",2014,6.3,"Chemnitz"
"Y_GE15","DED5",2014,8.3,"Leipzig"
"Y_GE15","DEE",2014,8.8,"Sachsen-Anhalt"
"Y_GE15","DEE0",2014,8.8,"Sachsen-Anhalt"
"Y_GE15","DEF",2014,4.6,"Schleswig-Holstein"
"Y_GE15","DEF0",2014,4.6,"Schleswig-Holstein"
"Y_GE15","DEG",2014,6,"Thüringen"
"Y_GE15","DEG0",2014,6,"Thüringen"
"Y_GE15","DK",2014,6.6,"Denmark"
"Y_GE15","DK0",2014,6.6,"Danmark"
"Y_GE15","DK01",2014,7.1,"Hovedstaden"
"Y_GE15","DK02",2014,6.3,"Sjælland"
"Y_GE15","DK03",2014,6.7,"Syddanmark"
"Y_GE15","DK04",2014,6.1,"Midtjylland"
"Y_GE15","DK05",2014,6.4,"Nordjylland"
"Y_GE15","EA17",2014,11.6,"Euro area (17 countries)"
"Y_GE15","EA18",2014,11.6,"Euro area (18 countries)"
"Y_GE15","EA19",2014,11.6,"Euro area (19 countries)"
"Y_GE15","EE",2014,7.4,"Estonia"
"Y_GE15","EE0",2014,7.4,"Eesti"
"Y_GE15","EE00",2014,7.4,"Eesti"
"Y_GE15","EL",2014,26.5,"Greece"
"Y_GE15","EL3",2014,27.3,"Attiki"
"Y_GE15","EL30",2014,27.3,"Attiki"
"Y_GE15","EL4",2014,22.5,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2014,22.3,"Voreio Aigaio"
"Y_GE15","EL42",2014,20.1,"Notio Aigaio"
"Y_GE15","EL43",2014,24,"Kriti"
"Y_GE15","EL5",2014,27.5,"Voreia Ellada"
"Y_GE15","EL51",2014,24.2,"Anatoliki Makedonia, Thraki"
"Y_GE15","EL52",2014,28.7,"Kentriki Makedonia"
"Y_GE15","EL53",2014,27.6,"Dytiki Makedonia"
"Y_GE15","EL54",2014,26.8,"Ipeiros"
"Y_GE15","EL6",2014,25.7,"Kentriki Ellada"
"Y_GE15","EL61",2014,25.4,"Thessalia"
"Y_GE15","EL62",2014,21.4,"Ionia Nisia"
"Y_GE15","EL63",2014,28.7,"Dytiki Ellada"
"Y_GE15","EL64",2014,26.8,"Sterea Ellada"
"Y_GE15","EL65",2014,23.4,"Peloponnisos"
"Y_GE15","ES",2014,24.4,"Spain"
"Y_GE15","ES1",2014,21.2,"Noroeste (ES)"
"Y_GE15","ES11",2014,21.7,"Galicia"
"Y_GE15","ES12",2014,21.1,"Principado de Asturias"
"Y_GE15","ES13",2014,19.4,"Cantabria"
"Y_GE15","ES2",2014,17.5,"Noreste (ES)"
"Y_GE15","ES21",2014,16.3,"País Vasco"
"Y_GE15","ES22",2014,15.7,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2014,18.2,"La Rioja"
"Y_GE15","ES24",2014,20.2,"Aragón"
"Y_GE15","ES3",2014,18.7,"Comunidad de Madrid"
"Y_GE15","ES30",2014,18.7,"Comunidad de Madrid"
"Y_GE15","ES4",2014,25.6,"Centro (ES)"
"Y_GE15","ES41",2014,20.8,"Castilla y León"
"Y_GE15","ES42",2014,29,"Castilla-la Mancha"
"Y_GE15","ES43",2014,29.8,"Extremadura"
"Y_GE15","ES5",2014,22.2,"Este (ES)"
"Y_GE15","ES51",2014,20.3,"Cataluña"
"Y_GE15","ES52",2014,25.8,"Comunidad Valenciana"
"Y_GE15","ES53",2014,20,"Illes Balears"
"Y_GE15","ES6",2014,33.5,"Sur (ES)"
"Y_GE15","ES61",2014,34.8,"Andalucía"
"Y_GE15","ES62",2014,26.6,"Región de Murcia"
"Y_GE15","ES63",2014,31.9,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2014,28.4,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2014,32.4,"Canarias (ES)"
"Y_GE15","ES70",2014,32.4,"Canarias (ES)"
"Y_GE15","EU15",2014,10.5,"European Union (15 countries)"
"Y_GE15","EU27",2014,10.2,"European Union (27 countries)"
"Y_GE15","EU28",2014,10.2,"European Union (28 countries)"
"Y_GE15","FI",2014,8.7,"Finland"
"Y_GE15","FI1",2014,8.7,"Manner-Suomi"
"Y_GE15","FI19",2014,8.7,"Länsi-Suomi"
"Y_GE15","FI1B",2014,7.3,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2014,9.4,"Etelä-Suomi"
"Y_GE15","FI1D",2014,10,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2014,NA,"Åland"
"Y_GE15","FI20",2014,NA,"Åland"
"Y_GE15","FR",2014,10.3,"France"
"Y_GE15","FR1",2014,9.7,"Île de France"
"Y_GE15","FR10",2014,9.7,"Île de France"
"Y_GE15","FR2",2014,10.5,"Bassin Parisien"
"Y_GE15","FR21",2014,11.4,"Champagne-Ardenne"
"Y_GE15","FR22",2014,11.6,"Picardie"
"Y_GE15","FR23",2014,11.9,"Haute-Normandie"
"Y_GE15","FR24",2014,9.5,"Centre (FR)"
"Y_GE15","FR25",2014,8.2,"Basse-Normandie"
"Y_GE15","FR26",2014,10.7,"Bourgogne"
"Y_GE15","FR3",2014,13.8,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2014,13.8,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2014,10.8,"Est (FR)"
"Y_GE15","FR41",2014,11.8,"Lorraine"
"Y_GE15","FR42",2014,10.1,"Alsace"
"Y_GE15","FR43",2014,9.8,"Franche-Comté"
"Y_GE15","FR5",2014,8.6,"Ouest (FR)"
"Y_GE15","FR51",2014,8.6,"Pays de la Loire"
"Y_GE15","FR52",2014,7.4,"Bretagne"
"Y_GE15","FR53",2014,10.9,"Poitou-Charentes"
"Y_GE15","FR6",2014,9.1,"Sud-Ouest (FR)"
"Y_GE15","FR61",2014,9,"Aquitaine"
"Y_GE15","FR62",2014,9.1,"Midi-Pyrénées"
"Y_GE15","FR63",2014,9.3,"Limousin"
"Y_GE15","FR7",2014,8.5,"Centre-Est (FR)"
"Y_GE15","FR71",2014,8.8,"Rhône-Alpes"
"Y_GE15","FR72",2014,7.4,"Auvergne"
"Y_GE15","FR8",2014,10.8,"Méditerranée"
"Y_GE15","FR81",2014,12.3,"Languedoc-Roussillon"
"Y_GE15","FR82",2014,10.1,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2014,9.9,"Corse"
"Y_GE15","FRA",2014,23.6,"Départements d'outre-mer"
"Y_GE15","FRA1",2014,23.9,"Guadeloupe"
"Y_GE15","FRA2",2014,19.4,"Martinique"
"Y_GE15","FRA3",2014,22.2,"Guyane"
"Y_GE15","FRA4",2014,26.4,"La Réunion"
"Y_GE15","FRA5",2014,19.6,"Mayotte"
"Y_GE15","HR",2014,17.3,"Croatia"
"Y_GE15","HR0",2014,17.3,"Hrvatska"
"Y_GE15","HR03",2014,17.2,"Jadranska Hrvatska"
"Y_GE15","HR04",2014,17.3,"Kontinentalna Hrvatska"
"Y_GE15","HU",2014,7.7,"Hungary"
"Y_GE15","HU1",2014,6.2,"Közép-Magyarország"
"Y_GE15","HU10",2014,6.2,"Közép-Magyarország"
"Y_GE15","HU2",2014,5.9,"Dunántúl"
"Y_GE15","HU21",2014,5.6,"Közép-Dunántúl"
"Y_GE15","HU22",2014,4.6,"Nyugat-Dunántúl"
"Y_GE15","HU23",2014,7.8,"Dél-Dunántúl"
"Y_GE15","HU3",2014,10.5,"Alföld és Észak"
"Y_GE15","HU31",2014,10.4,"Észak-Magyarország"
"Y_GE15","HU32",2014,11.8,"Észak-Alföld"
"Y_GE15","HU33",2014,9,"Dél-Alföld"
"Y_GE15","IE",2014,11.3,"Ireland"
"Y_GE15","IE0",2014,11.3,"Éire/Ireland"
"Y_GE15","IE01",2014,12.3,"Border, Midland and Western"
"Y_GE15","IE02",2014,10.9,"Southern and Eastern"
"Y_GE15","IS",2014,4.9,"Iceland"
"Y_GE15","IS0",2014,4.9,"Ísland"
"Y_GE15","IS00",2014,4.9,"Ísland"
"Y_GE15","IT",2014,12.7,"Italy"
"Y_GE15","ITC",2014,9.3,"Nord-Ovest"
"Y_GE15","ITC1",2014,11.3,"Piemonte"
"Y_GE15","ITC2",2014,8.9,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2014,10.8,"Liguria"
"Y_GE15","ITC4",2014,8.2,"Lombardia"
"Y_GE15","ITF",2014,20.4,"Sud"
"Y_GE15","ITF1",2014,12.6,"Abruzzo"
"Y_GE15","ITF2",2014,15.2,"Molise"
"Y_GE15","ITF3",2014,21.7,"Campania"
"Y_GE15","ITF4",2014,21.5,"Puglia"
"Y_GE15","ITF5",2014,14.7,"Basilicata"
"Y_GE15","ITF6",2014,23.4,"Calabria"
"Y_GE15","ITG",2014,21.2,"Isole"
"Y_GE15","ITG1",2014,22.2,"Sicilia"
"Y_GE15","ITG2",2014,18.6,"Sardegna"
"Y_GE15","ITH",2014,7.7,"Nord-Est"
"Y_GE15","ITH1",2014,4.4,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2014,6.9,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2014,7.5,"Veneto"
"Y_GE15","ITH4",2014,8,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2014,8.3,"Emilia-Romagna"
"Y_GE15","ITI",2014,11.4,"Centro (IT)"
"Y_GE15","ITI1",2014,10.1,"Toscana"
"Y_GE15","ITI2",2014,11.3,"Umbria"
"Y_GE15","ITI3",2014,10.1,"Marche"
"Y_GE15","ITI4",2014,12.5,"Lazio"
"Y_GE15","LT",2014,10.7,"Lithuania"
"Y_GE15","LT0",2014,10.7,"Lietuva"
"Y_GE15","LT00",2014,10.7,"Lietuva"
"Y_GE15","LU",2014,5.9,"Luxembourg"
"Y_GE15","LU0",2014,5.9,"Luxembourg"
"Y_GE15","LU00",2014,5.9,"Luxembourg"
"Y_GE15","LV",2014,10.8,"Latvia"
"Y_GE15","LV0",2014,10.8,"Latvija"
"Y_GE15","LV00",2014,10.8,"Latvija"
"Y_GE15","MK",2014,28,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2014,28,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2014,28,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2014,5.8,"Malta"
"Y_GE15","MT0",2014,5.8,"Malta"
"Y_GE15","MT00",2014,5.8,"Malta"
"Y_GE15","NL",2014,7.4,"Netherlands"
"Y_GE15","NL1",2014,8,"Noord-Nederland"
"Y_GE15","NL11",2014,8.6,"Groningen"
"Y_GE15","NL12",2014,7.9,"Friesland (NL)"
"Y_GE15","NL13",2014,7.3,"Drenthe"
"Y_GE15","NL2",2014,7.5,"Oost-Nederland"
"Y_GE15","NL21",2014,7.3,"Overijssel"
"Y_GE15","NL22",2014,6.9,"Gelderland"
"Y_GE15","NL23",2014,11,"Flevoland"
"Y_GE15","NL3",2014,7.4,"West-Nederland"
"Y_GE15","NL31",2014,6.4,"Utrecht"
"Y_GE15","NL32",2014,6.9,"Noord-Holland"
"Y_GE15","NL33",2014,8.4,"Zuid-Holland"
"Y_GE15","NL34",2014,5.4,"Zeeland"
"Y_GE15","NL4",2014,7.1,"Zuid-Nederland"
"Y_GE15","NL41",2014,7,"Noord-Brabant"
"Y_GE15","NL42",2014,7.4,"Limburg (NL)"
"Y_GE15","NO",2014,3.5,"Norway"
"Y_GE15","NO0",2014,3.5,"Norge"
"Y_GE15","NO01",2014,3.8,"Oslo og Akershus"
"Y_GE15","NO02",2014,2.9,"Hedmark og Oppland"
"Y_GE15","NO03",2014,4.1,"Sør-Østlandet"
"Y_GE15","NO04",2014,3.1,"Agder og Rogaland"
"Y_GE15","NO05",2014,3,"Vestlandet"
"Y_GE15","NO06",2014,3.8,"Trøndelag"
"Y_GE15","NO07",2014,3.3,"Nord-Norge"
"Y_GE15","PL",2014,9,"Poland"
"Y_GE15","PL1",2014,7.7,"Region Centralny"
"Y_GE15","PL11",2014,8.9,"Lódzkie"
"Y_GE15","PL12",2014,7.2,"Mazowieckie"
"Y_GE15","PL2",2014,8.8,"Region Poludniowy"
"Y_GE15","PL21",2014,9.1,"Malopolskie"
"Y_GE15","PL22",2014,8.6,"Slaskie"
"Y_GE15","PL3",2014,11.2,"Region Wschodni"
"Y_GE15","PL31",2014,9.9,"Lubelskie"
"Y_GE15","PL32",2014,14,"Podkarpackie"
"Y_GE15","PL33",2014,11.4,"Swietokrzyskie"
"Y_GE15","PL34",2014,9.1,"Podlaskie"
"Y_GE15","PL4",2014,8,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2014,7.7,"Wielkopolskie"
"Y_GE15","PL42",2014,8.4,"Zachodniopomorskie"
"Y_GE15","PL43",2014,8.3,"Lubuskie"
"Y_GE15","PL5",2014,8.8,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2014,9.1,"Dolnoslaskie"
"Y_GE15","PL52",2014,7.8,"Opolskie"
"Y_GE15","PL6",2014,9.6,"Region Pólnocny"
"Y_GE15","PL61",2014,10.7,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2014,9.8,"Warminsko-Mazurskie"
"Y_GE15","PL63",2014,8.6,"Pomorskie"
"Y_GE15","PT",2014,13.9,"Portugal"
"Y_GE15","PT1",2014,13.8,"Continente"
"Y_GE15","PT11",2014,14.8,"Norte"
"Y_GE15","PT15",2014,14.5,"Algarve"
"Y_GE15","PT16",2014,10.6,"Centro (PT)"
"Y_GE15","PT17",2014,14.9,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2014,14.3,"Alentejo"
"Y_GE15","PT2",2014,16.3,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2014,16.3,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2014,15,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2014,15,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2014,6.8,"Romania"
"Y_GE15","RO1",2014,6.2,"Macroregiunea unu"
"Y_GE15","RO11",2014,3.8,"Nord-Vest"
"Y_GE15","RO12",2014,9.2,"Centru"
"Y_GE15","RO2",2014,6.6,"Macroregiunea doi"
"Y_GE15","RO21",2014,4.2,"Nord-Est"
"Y_GE15","RO22",2014,10.4,"Sud-Est"
"Y_GE15","RO3",2014,8.2,"Macroregiunea trei"
"Y_GE15","RO31",2014,9,"Sud - Muntenia"
"Y_GE15","RO32",2014,7.2,"Bucuresti - Ilfov"
"Y_GE15","RO4",2014,5.7,"Macroregiunea patru"
"Y_GE15","RO41",2014,6.5,"Sud-Vest Oltenia"
"Y_GE15","RO42",2014,4.8,"Vest"
"Y_GE15","SE",2014,8,"Sweden"
"Y_GE15","SE1",2014,7.6,"Östra Sverige"
"Y_GE15","SE11",2014,7.1,"Stockholm"
"Y_GE15","SE12",2014,8.3,"Östra Mellansverige"
"Y_GE15","SE2",2014,8.3,"Södra Sverige"
"Y_GE15","SE21",2014,6.7,"Småland med öarna"
"Y_GE15","SE22",2014,10,"Sydsverige"
"Y_GE15","SE23",2014,7.6,"Västsverige"
"Y_GE15","SE3",2014,8,"Norra Sverige"
"Y_GE15","SE31",2014,8.6,"Norra Mellansverige"
"Y_GE15","SE32",2014,7.4,"Mellersta Norrland"
"Y_GE15","SE33",2014,7.4,"Övre Norrland"
"Y_GE15","SI",2014,9.7,"Slovenia"
"Y_GE15","SI0",2014,9.7,"Slovenija"
"Y_GE15","SI03",2014,11,"Vzhodna Slovenija"
"Y_GE15","SI04",2014,8.1,"Zahodna Slovenija"
"Y_GE15","SK",2014,13.2,"Slovakia"
"Y_GE15","SK0",2014,13.2,"Slovensko"
"Y_GE15","SK01",2014,6,"Bratislavský kraj"
"Y_GE15","SK02",2014,11,"Západné Slovensko"
"Y_GE15","SK03",2014,15.9,"Stredné Slovensko"
"Y_GE15","SK04",2014,16.6,"Východné Slovensko"
"Y_GE15","TR",2014,9.9,"Turkey"
"Y_GE15","TR1",2014,11.9,"Istanbul"
"Y_GE15","TR10",2014,11.9,"Istanbul"
"Y_GE15","TR2",2014,6.7,"Bati Marmara"
"Y_GE15","TR21",2014,7.6,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2014,5.6,"Balikesir, Çanakkale"
"Y_GE15","TR3",2014,9,"Ege"
"Y_GE15","TR31",2014,13.8,"Izmir"
"Y_GE15","TR32",2014,7.2,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2014,3.9,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2014,8,"Dogu Marmara"
"Y_GE15","TR41",2014,6.2,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2014,9.9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2014,9.8,"Bati Anadolu"
"Y_GE15","TR51",2014,11.5,"Ankara"
"Y_GE15","TR52",2014,5.5,"Konya, Karaman"
"Y_GE15","TR6",2014,11.1,"Akdeniz"
"Y_GE15","TR61",2014,8.4,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2014,10.7,"Adana, Mersin"
"Y_GE15","TR63",2014,15.3,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2014,8.8,"Orta Anadolu"
"Y_GE15","TR71",2014,7.6,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2014,9.5,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2014,6.2,"Bati Karadeniz"
"Y_GE15","TR81",2014,6,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2014,6.5,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2014,6.2,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2014,6.2,"Dogu Karadeniz"
"Y_GE15","TR90",2014,6.2,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2014,5.2,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2014,7.3,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2014,3.3,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2014,10.6,"Ortadogu Anadolu"
"Y_GE15","TRB1",2014,7.5,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2014,13.4,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2014,15.6,"Güneydogu Anadolu"
"Y_GE15","TRC1",2014,8.1,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2014,17.5,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2014,24,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2014,6.1,"United Kingdom"
"Y_GE15","UKC",2014,9,"North East (UK)"
"Y_GE15","UKC1",2014,9.8,"Tees Valley and Durham"
"Y_GE15","UKC2",2014,8.3,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2014,6.7,"North West (UK)"
"Y_GE15","UKD1",2014,5,"Cumbria"
"Y_GE15","UKD3",2014,7.9,"Greater Manchester"
"Y_GE15","UKD4",2014,6.5,"Lancashire"
"Y_GE15","UKD6",2014,3.4,"Cheshire"
"Y_GE15","UKD7",2014,7.4,"Merseyside"
"Y_GE15","UKE",2014,7.2,"Yorkshire and The Humber"
"Y_GE15","UKE1",2014,8,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2014,4.6,"North Yorkshire"
"Y_GE15","UKE3",2014,8.8,"South Yorkshire"
"Y_GE15","UKE4",2014,6.7,"West Yorkshire"
"Y_GE15","UKF",2014,5.5,"East Midlands (UK)"
"Y_GE15","UKF1",2014,6.1,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2014,5.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2014,4.6,"Lincolnshire"
"Y_GE15","UKG",2014,7.2,"West Midlands (UK)"
"Y_GE15","UKG1",2014,4.4,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2014,5.3,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2014,9.7,"West Midlands"
"Y_GE15","UKH",2014,5.1,"East of England"
"Y_GE15","UKH1",2014,5,"East Anglia"
"Y_GE15","UKH2",2014,4.3,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2014,6.2,"Essex"
"Y_GE15","UKI",2014,6.8,"London"
"Y_GE15","UKI3",2014,6.2,"Inner London - West"
"Y_GE15","UKI4",2014,7.8,"Inner London - East"
"Y_GE15","UKI5",2014,7.4,"Outer London - East and North East"
"Y_GE15","UKI6",2014,5.9,"Outer London - South"
"Y_GE15","UKI7",2014,6.2,"Outer London - West and North West"
"Y_GE15","UKJ",2014,4.6,"South East (UK)"
"Y_GE15","UKJ1",2014,4.2,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2014,4.6,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2014,4.2,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2014,5.7,"Kent"
"Y_GE15","UKK",2014,4.7,"South West (UK)"
"Y_GE15","UKK1",2014,4.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2014,4.5,"Dorset and Somerset"
"Y_GE15","UKK3",2014,3.8,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2014,5,"Devon"
"Y_GE15","UKL",2014,6.6,"Wales"
"Y_GE15","UKL1",2014,6.9,"West Wales and The Valleys"
"Y_GE15","UKL2",2014,6.1,"East Wales"
"Y_GE15","UKM",2014,5.9,"Scotland"
"Y_GE15","UKM2",2014,5.6,"Eastern Scotland"
"Y_GE15","UKM3",2014,7.1,"South Western Scotland"
"Y_GE15","UKM5",2014,4,"North Eastern Scotland"
"Y_GE15","UKM6",2014,4.4,"Highlands and Islands"
"Y_GE15","UKN",2014,6.4,"Northern Ireland (UK)"
"Y_GE15","UKN0",2014,6.4,"Northern Ireland (UK)"
"Y_GE25","AT",2014,4.9,"Austria"
"Y_GE25","AT1",2014,6.5,"Ostösterreich"
"Y_GE25","AT11",2014,4.1,"Burgenland (AT)"
"Y_GE25","AT12",2014,4.2,"Niederösterreich"
"Y_GE25","AT13",2014,9.1,"Wien"
"Y_GE25","AT2",2014,4.8,"Südösterreich"
"Y_GE25","AT21",2014,5.4,"Kärnten"
"Y_GE25","AT22",2014,4.5,"Steiermark"
"Y_GE25","AT3",2014,3.1,"Westösterreich"
"Y_GE25","AT31",2014,3.4,"Oberösterreich"
"Y_GE25","AT32",2014,3.2,"Salzburg"
"Y_GE25","AT33",2014,2.8,"Tirol"
"Y_GE25","AT34",2014,2.5,"Vorarlberg"
"Y_GE25","BE",2014,7.2,"Belgium"
"Y_GE25","BE1",2014,16.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2014,16.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2014,4.1,"Vlaams Gewest"
"Y_GE25","BE21",2014,5.1,"Prov. Antwerpen"
"Y_GE25","BE22",2014,4.7,"Prov. Limburg (BE)"
"Y_GE25","BE23",2014,3.2,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2014,4,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2014,3.2,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2014,10,"Région wallonne"
"Y_GE25","BE31",2014,7.8,"Prov. Brabant Wallon"
"Y_GE25","BE32",2014,12.3,"Prov. Hainaut"
"Y_GE25","BE33",2014,10.5,"Prov. Liège"
"Y_GE25","BE34",2014,7,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2014,7,"Prov. Namur"
"Y_GE25","BG",2014,10.6,"Bulgaria"
"Y_GE25","BG3",2014,12.1,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2014,13.3,"Severozapaden"
"Y_GE25","BG32",2014,12.5,"Severen tsentralen"
"Y_GE25","BG33",2014,12,"Severoiztochen"
"Y_GE25","BG34",2014,10.9,"Yugoiztochen"
"Y_GE25","BG4",2014,9.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2014,8.4,"Yugozapaden"
"Y_GE25","BG42",2014,10.8,"Yuzhen tsentralen"
"Y_GE25","CH",2014,3.9,"Switzerland"
"Y_GE25","CH0",2014,3.9,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2014,5.6,"Région lémanique"
"Y_GE25","CH02",2014,3.6,"Espace Mittelland"
"Y_GE25","CH03",2014,3.9,"Nordwestschweiz"
"Y_GE25","CH04",2014,3.8,"Zürich"
"Y_GE25","CH05",2014,2.8,"Ostschweiz"
"Y_GE25","CH06",2014,2.9,"Zentralschweiz"
"Y_GE25","CH07",2014,5.6,"Ticino"
"Y_GE25","CY",2014,13.9,"Cyprus"
"Y_GE25","CY0",2014,13.9,"Kypros"
"Y_GE25","CY00",2014,13.9,"Kypros"
"Y_GE25","CZ",2014,5.4,"Czech Republic"
"Y_GE25","CZ0",2014,5.4,"Ceská republika"
"Y_GE25","CZ01",2014,2.1,"Praha"
"Y_GE25","CZ02",2014,4.6,"Strední Cechy"
"Y_GE25","CZ03",2014,4.8,"Jihozápad"
"Y_GE25","CZ04",2014,7.6,"Severozápad"
"Y_GE25","CZ05",2014,5.5,"Severovýchod"
"Y_GE25","CZ06",2014,5.3,"Jihovýchod"
"Y_GE25","CZ07",2014,6.3,"Strední Morava"
"Y_GE25","CZ08",2014,7.8,"Moravskoslezsko"
"Y_GE25","DE",2014,4.7,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2014,2.9,"Baden-Württemberg"
"Y_GE25","DE11",2014,2.9,"Stuttgart"
"Y_GE25","DE12",2014,3.3,"Karlsruhe"
"Y_GE25","DE13",2014,2.7,"Freiburg"
"Y_GE25","DE14",2014,2.2,"Tübingen"
"Y_GE25","DE2",2014,2.7,"Bayern"
"Y_GE25","DE21",2014,2.4,"Oberbayern"
"Y_GE25","DE22",2014,2.7,"Niederbayern"
"Y_GE25","DE23",2014,2.6,"Oberpfalz"
"Y_GE25","DE24",2014,3.7,"Oberfranken"
"Y_GE25","DE25",2014,2.8,"Mittelfranken"
"Y_GE25","DE26",2014,2.7,"Unterfranken"
"Y_GE25","DE27",2014,2.8,"Schwaben"
"Y_GE25","DE3",2014,9.3,"Berlin"
"Y_GE25","DE30",2014,9.3,"Berlin"
"Y_GE25","DE4",2014,6.4,"Brandenburg"
"Y_GE25","DE40",2014,6.4,"Brandenburg"
"Y_GE25","DE5",2014,6,"Bremen"
"Y_GE25","DE50",2014,6,"Bremen"
"Y_GE25","DE6",2014,4.7,"Hamburg"
"Y_GE25","DE60",2014,4.7,"Hamburg"
"Y_GE25","DE7",2014,3.9,"Hessen"
"Y_GE25","DE71",2014,3.9,"Darmstadt"
"Y_GE25","DE72",2014,3.6,"Gießen"
"Y_GE25","DE73",2014,3.9,"Kassel"
"Y_GE25","DE8",2014,9.4,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2014,9.4,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2014,4.4,"Niedersachsen"
"Y_GE25","DE91",2014,5.3,"Braunschweig"
"Y_GE25","DE92",2014,4.9,"Hannover"
"Y_GE25","DE93",2014,3.7,"Lüneburg"
"Y_GE25","DE94",2014,3.8,"Weser-Ems"
"Y_GE25","DEA",2014,5.2,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2014,6.1,"Düsseldorf"
"Y_GE25","DEA2",2014,4.8,"Köln"
"Y_GE25","DEA3",2014,4.3,"Münster"
"Y_GE25","DEA4",2014,4.5,"Detmold"
"Y_GE25","DEA5",2014,5.2,"Arnsberg"
"Y_GE25","DEB",2014,3.4,"Rheinland-Pfalz"
"Y_GE25","DEB1",2014,3.5,"Koblenz"
"Y_GE25","DEB2",2014,2.5,"Trier"
"Y_GE25","DEB3",2014,3.5,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2014,5.5,"Saarland"
"Y_GE25","DEC0",2014,5.5,"Saarland"
"Y_GE25","DED",2014,6.9,"Sachsen"
"Y_GE25","DED2",2014,6.9,"Dresden"
"Y_GE25","DED4",2014,6.2,"Chemnitz"
"Y_GE25","DED5",2014,8,"Leipzig"
"Y_GE25","DEE",2014,8.5,"Sachsen-Anhalt"
"Y_GE25","DEE0",2014,8.5,"Sachsen-Anhalt"
"Y_GE25","DEF",2014,4.1,"Schleswig-Holstein"
"Y_GE25","DEF0",2014,4.1,"Schleswig-Holstein"
"Y_GE25","DEG",2014,5.8,"Thüringen"
"Y_GE25","DEG0",2014,5.8,"Thüringen"
"Y_GE25","DK",2014,5.5,"Denmark"
"Y_GE25","DK0",2014,5.5,"Danmark"
"Y_GE25","DK01",2014,6.1,"Hovedstaden"
"Y_GE25","DK02",2014,5,"Sjælland"
"Y_GE25","DK03",2014,5.6,"Syddanmark"
"Y_GE25","DK04",2014,5,"Midtjylland"
"Y_GE25","DK05",2014,5.1,"Nordjylland"
"Y_GE25","EA17",2014,10.4,"Euro area (17 countries)"
"Y_GE25","EA18",2014,10.4,"Euro area (18 countries)"
"Y_GE25","EA19",2014,10.4,"Euro area (19 countries)"
"Y_GE25","EE",2014,6.7,"Estonia"
"Y_GE25","EE0",2014,6.7,"Eesti"
"Y_GE25","EE00",2014,6.7,"Eesti"
"Y_GE25","EL",2014,24.7,"Greece"
"Y_GE25","EL3",2014,25.7,"Attiki"
"Y_GE25","EL30",2014,25.7,"Attiki"
"Y_GE25","EL4",2014,21.2,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2014,20.8,"Voreio Aigaio"
"Y_GE25","EL42",2014,19.6,"Notio Aigaio"
"Y_GE25","EL43",2014,22.2,"Kriti"
"Y_GE25","EL5",2014,25.8,"Voreia Ellada"
"Y_GE25","EL51",2014,22,"Anatoliki Makedonia, Thraki"
"Y_GE25","EL52",2014,27.2,"Kentriki Makedonia"
"Y_GE25","EL53",2014,26.3,"Dytiki Makedonia"
"Y_GE25","EL54",2014,24.2,"Ipeiros"
"Y_GE25","EL6",2014,23.5,"Kentriki Ellada"
"Y_GE25","EL61",2014,23.3,"Thessalia"
"Y_GE25","EL62",2014,19.6,"Ionia Nisia"
"Y_GE25","EL63",2014,26,"Dytiki Ellada"
"Y_GE25","EL64",2014,24.3,"Sterea Ellada"
"Y_GE25","EL65",2014,21.5,"Peloponnisos"
"Y_GE25","ES",2014,22.3,"Spain"
"Y_GE25","ES1",2014,19.8,"Noroeste (ES)"
"Y_GE25","ES11",2014,20.1,"Galicia"
"Y_GE25","ES12",2014,20,"Principado de Asturias"
"Y_GE25","ES13",2014,18,"Cantabria"
"Y_GE25","ES2",2014,15.8,"Noreste (ES)"
"Y_GE25","ES21",2014,15,"País Vasco"
"Y_GE25","ES22",2014,13.8,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2014,16.3,"La Rioja"
"Y_GE25","ES24",2014,18,"Aragón"
"Y_GE25","ES3",2014,16.7,"Comunidad de Madrid"
"Y_GE25","ES30",2014,16.7,"Comunidad de Madrid"
"Y_GE25","ES4",2014,23.2,"Centro (ES)"
"Y_GE25","ES41",2014,19,"Castilla y León"
"Y_GE25","ES42",2014,26.1,"Castilla-la Mancha"
"Y_GE25","ES43",2014,27.5,"Extremadura"
"Y_GE25","ES5",2014,20,"Este (ES)"
"Y_GE25","ES51",2014,18.2,"Cataluña"
"Y_GE25","ES52",2014,23.4,"Comunidad Valenciana"
"Y_GE25","ES53",2014,18.1,"Illes Balears"
"Y_GE25","ES6",2014,31.1,"Sur (ES)"
"Y_GE25","ES61",2014,32.4,"Andalucía"
"Y_GE25","ES62",2014,24.4,"Región de Murcia"
"Y_GE25","ES63",2014,28.2,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2014,26.1,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2014,30.4,"Canarias (ES)"
"Y_GE25","ES70",2014,30.4,"Canarias (ES)"
"Y_GE25","EU15",2014,9.2,"European Union (15 countries)"
"Y_GE25","EU27",2014,8.9,"European Union (27 countries)"
"Y_GE25","EU28",2014,8.9,"European Union (28 countries)"
"Y_GE25","FI",2014,7,"Finland"
"Y_GE25","FI1",2014,7,"Manner-Suomi"
"Y_GE25","FI19",2014,7,"Länsi-Suomi"
"Y_GE25","FI1B",2014,5.8,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2014,7.6,"Etelä-Suomi"
"Y_GE25","FI1D",2014,8.2,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2014,NA,"Åland"
"Y_GE25","FI20",2014,NA,"Åland"
"Y_GE25","FR",2014,8.9,"France"
"Y_GE25","FR1",2014,8.7,"Île de France"
"Y_GE25","FR10",2014,8.7,"Île de France"
"Y_GE25","FR2",2014,8.9,"Bassin Parisien"
"Y_GE25","FR21",2014,9.6,"Champagne-Ardenne"
"Y_GE25","FR22",2014,9.7,"Picardie"
"Y_GE25","FR23",2014,10.3,"Haute-Normandie"
"Y_GE25","FR24",2014,8.2,"Centre (FR)"
"Y_GE25","FR25",2014,6.6,"Basse-Normandie"
"Y_GE25","FR26",2014,9.2,"Bourgogne"
"Y_GE25","FR3",2014,11.9,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2014,11.9,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2014,9.1,"Est (FR)"
"Y_GE25","FR41",2014,10.3,"Lorraine"
"Y_GE25","FR42",2014,8.1,"Alsace"
"Y_GE25","FR43",2014,8.7,"Franche-Comté"
"Y_GE25","FR5",2014,7.2,"Ouest (FR)"
"Y_GE25","FR51",2014,7.2,"Pays de la Loire"
"Y_GE25","FR52",2014,6.2,"Bretagne"
"Y_GE25","FR53",2014,9,"Poitou-Charentes"
"Y_GE25","FR6",2014,7.8,"Sud-Ouest (FR)"
"Y_GE25","FR61",2014,7.6,"Aquitaine"
"Y_GE25","FR62",2014,7.9,"Midi-Pyrénées"
"Y_GE25","FR63",2014,7.4,"Limousin"
"Y_GE25","FR7",2014,7.3,"Centre-Est (FR)"
"Y_GE25","FR71",2014,7.5,"Rhône-Alpes"
"Y_GE25","FR72",2014,6.2,"Auvergne"
"Y_GE25","FR8",2014,9.3,"Méditerranée"
"Y_GE25","FR81",2014,10.5,"Languedoc-Roussillon"
"Y_GE25","FR82",2014,8.7,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2014,7.9,"Corse"
"Y_GE25","FRA",2014,20.5,"Départements d'outre-mer"
"Y_GE25","FRA1",2014,21.2,"Guadeloupe"
"Y_GE25","FRA2",2014,17,"Martinique"
"Y_GE25","FRA3",2014,19.8,"Guyane"
"Y_GE25","FRA4",2014,22.6,"La Réunion"
"Y_GE25","FRA5",2014,16.5,"Mayotte"
"Y_GE25","HR",2014,14.6,"Croatia"
"Y_GE25","HR0",2014,14.6,"Hrvatska"
"Y_GE25","HR03",2014,14.4,"Jadranska Hrvatska"
"Y_GE25","HR04",2014,14.7,"Kontinentalna Hrvatska"
"Y_GE25","HU",2014,6.7,"Hungary"
"Y_GE25","HU1",2014,5.6,"Közép-Magyarország"
"Y_GE25","HU10",2014,5.6,"Közép-Magyarország"
"Y_GE25","HU2",2014,5.1,"Dunántúl"
"Y_GE25","HU21",2014,4.7,"Közép-Dunántúl"
"Y_GE25","HU22",2014,3.9,"Nyugat-Dunántúl"
"Y_GE25","HU23",2014,6.9,"Dél-Dunántúl"
"Y_GE25","HU3",2014,9,"Alföld és Észak"
"Y_GE25","HU31",2014,9.1,"Észak-Magyarország"
"Y_GE25","HU32",2014,10.1,"Észak-Alföld"
"Y_GE25","HU33",2014,7.6,"Dél-Alföld"
"Y_GE25","IE",2014,10,"Ireland"
"Y_GE25","IE0",2014,10,"Éire/Ireland"
"Y_GE25","IE01",2014,10.6,"Border, Midland and Western"
"Y_GE25","IE02",2014,9.8,"Southern and Eastern"
"Y_GE25","IS",2014,3.9,"Iceland"
"Y_GE25","IS0",2014,3.9,"Ísland"
"Y_GE25","IS00",2014,3.9,"Ísland"
"Y_GE25","IT",2014,10.6,"Italy"
"Y_GE25","ITC",2014,7.6,"Nord-Ovest"
"Y_GE25","ITC1",2014,9.3,"Piemonte"
"Y_GE25","ITC2",2014,7.4,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2014,9,"Liguria"
"Y_GE25","ITC4",2014,6.7,"Lombardia"
"Y_GE25","ITF",2014,17.4,"Sud"
"Y_GE25","ITF1",2014,10.5,"Abruzzo"
"Y_GE25","ITF2",2014,13.1,"Molise"
"Y_GE25","ITF3",2014,18.7,"Campania"
"Y_GE25","ITF4",2014,18.1,"Puglia"
"Y_GE25","ITF5",2014,12.6,"Basilicata"
"Y_GE25","ITF6",2014,20.2,"Calabria"
"Y_GE25","ITG",2014,18.3,"Isole"
"Y_GE25","ITG1",2014,19,"Sicilia"
"Y_GE25","ITG2",2014,16.4,"Sardegna"
"Y_GE25","ITH",2014,6.3,"Nord-Est"
"Y_GE25","ITH1",2014,3.6,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2014,5.5,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2014,6.1,"Veneto"
"Y_GE25","ITH4",2014,6.9,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2014,6.8,"Emilia-Romagna"
"Y_GE25","ITI",2014,9.6,"Centro (IT)"
"Y_GE25","ITI1",2014,8.5,"Toscana"
"Y_GE25","ITI2",2014,9.4,"Umbria"
"Y_GE25","ITI3",2014,8.5,"Marche"
"Y_GE25","ITI4",2014,10.5,"Lazio"
"Y_GE25","LT",2014,9.9,"Lithuania"
"Y_GE25","LT0",2014,9.9,"Lietuva"
"Y_GE25","LT00",2014,9.9,"Lietuva"
"Y_GE25","LU",2014,4.8,"Luxembourg"
"Y_GE25","LU0",2014,4.8,"Luxembourg"
"Y_GE25","LU00",2014,4.8,"Luxembourg"
"Y_GE25","LV",2014,10,"Latvia"
"Y_GE25","LV0",2014,10,"Latvija"
"Y_GE25","LV00",2014,10,"Latvija"
"Y_GE25","MK",2014,25.3,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2014,25.3,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2014,25.3,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2014,4.8,"Malta"
"Y_GE25","MT0",2014,4.8,"Malta"
"Y_GE25","MT00",2014,4.8,"Malta"
"Y_GE25","NL",2014,6.4,"Netherlands"
"Y_GE25","NL1",2014,6.8,"Noord-Nederland"
"Y_GE25","NL11",2014,7.2,"Groningen"
"Y_GE25","NL12",2014,6.9,"Friesland (NL)"
"Y_GE25","NL13",2014,6.2,"Drenthe"
"Y_GE25","NL2",2014,6.6,"Oost-Nederland"
"Y_GE25","NL21",2014,6.3,"Overijssel"
"Y_GE25","NL22",2014,6.3,"Gelderland"
"Y_GE25","NL23",2014,9.1,"Flevoland"
"Y_GE25","NL3",2014,6.4,"West-Nederland"
"Y_GE25","NL31",2014,5.4,"Utrecht"
"Y_GE25","NL32",2014,6,"Noord-Holland"
"Y_GE25","NL33",2014,7.3,"Zuid-Holland"
"Y_GE25","NL34",2014,4.7,"Zeeland"
"Y_GE25","NL4",2014,6.2,"Zuid-Nederland"
"Y_GE25","NL41",2014,6.2,"Noord-Brabant"
"Y_GE25","NL42",2014,6.2,"Limburg (NL)"
"Y_GE25","NO",2014,2.8,"Norway"
"Y_GE25","NO0",2014,2.8,"Norge"
"Y_GE25","NO01",2014,3.3,"Oslo og Akershus"
"Y_GE25","NO02",2014,2.3,"Hedmark og Oppland"
"Y_GE25","NO03",2014,3.3,"Sør-Østlandet"
"Y_GE25","NO04",2014,2.5,"Agder og Rogaland"
"Y_GE25","NO05",2014,2.3,"Vestlandet"
"Y_GE25","NO06",2014,3.2,"Trøndelag"
"Y_GE25","NO07",2014,2.2,"Nord-Norge"
"Y_GE25","PL",2014,7.6,"Poland"
"Y_GE25","PL1",2014,6.8,"Region Centralny"
"Y_GE25","PL11",2014,7.9,"Lódzkie"
"Y_GE25","PL12",2014,6.3,"Mazowieckie"
"Y_GE25","PL2",2014,7.4,"Region Poludniowy"
"Y_GE25","PL21",2014,7.5,"Malopolskie"
"Y_GE25","PL22",2014,7.4,"Slaskie"
"Y_GE25","PL3",2014,9.3,"Region Wschodni"
"Y_GE25","PL31",2014,8.1,"Lubelskie"
"Y_GE25","PL32",2014,11.5,"Podkarpackie"
"Y_GE25","PL33",2014,9.8,"Swietokrzyskie"
"Y_GE25","PL34",2014,7.7,"Podlaskie"
"Y_GE25","PL4",2014,6.6,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2014,6.3,"Wielkopolskie"
"Y_GE25","PL42",2014,7.2,"Zachodniopomorskie"
"Y_GE25","PL43",2014,6.9,"Lubuskie"
"Y_GE25","PL5",2014,7.7,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2014,8,"Dolnoslaskie"
"Y_GE25","PL52",2014,6.7,"Opolskie"
"Y_GE25","PL6",2014,8.2,"Region Pólnocny"
"Y_GE25","PL61",2014,9,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2014,8.5,"Warminsko-Mazurskie"
"Y_GE25","PL63",2014,7.3,"Pomorskie"
"Y_GE25","PT",2014,12.3,"Portugal"
"Y_GE25","PT1",2014,12.2,"Continente"
"Y_GE25","PT11",2014,13,"Norte"
"Y_GE25","PT15",2014,13.1,"Algarve"
"Y_GE25","PT16",2014,9.4,"Centro (PT)"
"Y_GE25","PT17",2014,13.4,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2014,12.7,"Alentejo"
"Y_GE25","PT2",2014,13.3,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2014,13.3,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2014,12.4,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2014,12.4,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2014,5.5,"Romania"
"Y_GE25","RO1",2014,4.8,"Macroregiunea unu"
"Y_GE25","RO11",2014,3,"Nord-Vest"
"Y_GE25","RO12",2014,7.1,"Centru"
"Y_GE25","RO2",2014,5.6,"Macroregiunea doi"
"Y_GE25","RO21",2014,3.4,"Nord-Est"
"Y_GE25","RO22",2014,8.8,"Sud-Est"
"Y_GE25","RO3",2014,6.6,"Macroregiunea trei"
"Y_GE25","RO31",2014,6.9,"Sud - Muntenia"
"Y_GE25","RO32",2014,6.2,"Bucuresti - Ilfov"
"Y_GE25","RO4",2014,4.5,"Macroregiunea patru"
"Y_GE25","RO41",2014,5.2,"Sud-Vest Oltenia"
"Y_GE25","RO42",2014,3.5,"Vest"
"Y_GE25","SE",2014,5.7,"Sweden"
"Y_GE25","SE1",2014,5.5,"Östra Sverige"
"Y_GE25","SE11",2014,5.3,"Stockholm"
"Y_GE25","SE12",2014,5.8,"Östra Mellansverige"
"Y_GE25","SE2",2014,6,"Södra Sverige"
"Y_GE25","SE21",2014,4.6,"Småland med öarna"
"Y_GE25","SE22",2014,7.6,"Sydsverige"
"Y_GE25","SE23",2014,5.4,"Västsverige"
"Y_GE25","SE3",2014,5.7,"Norra Sverige"
"Y_GE25","SE31",2014,6.2,"Norra Mellansverige"
"Y_GE25","SE32",2014,5.4,"Mellersta Norrland"
"Y_GE25","SE33",2014,5.1,"Övre Norrland"
"Y_GE25","SI",2014,8.9,"Slovenia"
"Y_GE25","SI0",2014,8.9,"Slovenija"
"Y_GE25","SI03",2014,10.1,"Vzhodna Slovenija"
"Y_GE25","SI04",2014,7.5,"Zahodna Slovenija"
"Y_GE25","SK",2014,11.8,"Slovakia"
"Y_GE25","SK0",2014,11.8,"Slovensko"
"Y_GE25","SK01",2014,5.5,"Bratislavský kraj"
"Y_GE25","SK02",2014,9.8,"Západné Slovensko"
"Y_GE25","SK03",2014,14.4,"Stredné Slovensko"
"Y_GE25","SK04",2014,14.9,"Východné Slovensko"
"Y_GE25","TR",2014,8.3,"Turkey"
"Y_GE25","TR1",2014,10.3,"Istanbul"
"Y_GE25","TR10",2014,10.3,"Istanbul"
"Y_GE25","TR2",2014,5.5,"Bati Marmara"
"Y_GE25","TR21",2014,6.7,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2014,4.3,"Balikesir, Çanakkale"
"Y_GE25","TR3",2014,7.7,"Ege"
"Y_GE25","TR31",2014,12.3,"Izmir"
"Y_GE25","TR32",2014,6,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2014,3,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2014,6.6,"Dogu Marmara"
"Y_GE25","TR41",2014,5.3,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2014,8,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2014,8.4,"Bati Anadolu"
"Y_GE25","TR51",2014,10,"Ankara"
"Y_GE25","TR52",2014,4.4,"Konya, Karaman"
"Y_GE25","TR6",2014,9.5,"Akdeniz"
"Y_GE25","TR61",2014,7.3,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2014,9.2,"Adana, Mersin"
"Y_GE25","TR63",2014,13.1,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2014,7.4,"Orta Anadolu"
"Y_GE25","TR71",2014,6.5,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2014,8,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2014,5,"Bati Karadeniz"
"Y_GE25","TR81",2014,4.5,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2014,5,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2014,5.2,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2014,4.7,"Dogu Karadeniz"
"Y_GE25","TR90",2014,4.7,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2014,4.2,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2014,5.9,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2014,2.6,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2014,8.4,"Ortadogu Anadolu"
"Y_GE25","TRB1",2014,6,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2014,10.8,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2014,13.4,"Güneydogu Anadolu"
"Y_GE25","TRC1",2014,5.9,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2014,16.6,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2014,20.3,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2014,4.4,"United Kingdom"
"Y_GE25","UKC",2014,6.4,"North East (UK)"
"Y_GE25","UKC1",2014,6.9,"Tees Valley and Durham"
"Y_GE25","UKC2",2014,5.9,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2014,5,"North West (UK)"
"Y_GE25","UKD1",2014,3.8,"Cumbria"
"Y_GE25","UKD3",2014,5.9,"Greater Manchester"
"Y_GE25","UKD4",2014,5.1,"Lancashire"
"Y_GE25","UKD6",2014,2.6,"Cheshire"
"Y_GE25","UKD7",2014,5.3,"Merseyside"
"Y_GE25","UKE",2014,5.3,"Yorkshire and The Humber"
"Y_GE25","UKE1",2014,6.2,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2014,3.3,"North Yorkshire"
"Y_GE25","UKE3",2014,6.5,"South Yorkshire"
"Y_GE25","UKE4",2014,4.9,"West Yorkshire"
"Y_GE25","UKF",2014,4.2,"East Midlands (UK)"
"Y_GE25","UKF1",2014,4.4,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2014,4.1,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2014,3.9,"Lincolnshire"
"Y_GE25","UKG",2014,5,"West Midlands (UK)"
"Y_GE25","UKG1",2014,2.9,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2014,4.1,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2014,6.6,"West Midlands"
"Y_GE25","UKH",2014,3.6,"East of England"
"Y_GE25","UKH1",2014,3.4,"East Anglia"
"Y_GE25","UKH2",2014,3,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2014,4.6,"Essex"
"Y_GE25","UKI",2014,5.3,"London"
"Y_GE25","UKI3",2014,5.6,"Inner London - West"
"Y_GE25","UKI4",2014,6.2,"Inner London - East"
"Y_GE25","UKI5",2014,5.5,"Outer London - East and North East"
"Y_GE25","UKI6",2014,4.2,"Outer London - South"
"Y_GE25","UKI7",2014,4.5,"Outer London - West and North West"
"Y_GE25","UKJ",2014,3.1,"South East (UK)"
"Y_GE25","UKJ1",2014,3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2014,3,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2014,2.8,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2014,3.9,"Kent"
"Y_GE25","UKK",2014,3.1,"South West (UK)"
"Y_GE25","UKK1",2014,3.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2014,2.6,"Dorset and Somerset"
"Y_GE25","UKK3",2014,2.7,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2014,3.1,"Devon"
"Y_GE25","UKL",2014,4.5,"Wales"
"Y_GE25","UKL1",2014,4.8,"West Wales and The Valleys"
"Y_GE25","UKL2",2014,4.1,"East Wales"
"Y_GE25","UKM",2014,4.1,"Scotland"
"Y_GE25","UKM2",2014,3.6,"Eastern Scotland"
"Y_GE25","UKM3",2014,5.1,"South Western Scotland"
"Y_GE25","UKM5",2014,3.6,"North Eastern Scotland"
"Y_GE25","UKM6",2014,2.7,"Highlands and Islands"
"Y_GE25","UKN",2014,4.5,"Northern Ireland (UK)"
"Y_GE25","UKN0",2014,4.5,"Northern Ireland (UK)"
"Y15-24","AT",2013,9.7,"Austria"
"Y15-24","AT1",2013,12.9,"Ostösterreich"
"Y15-24","AT11",2013,NA,"Burgenland (AT)"
"Y15-24","AT12",2013,10.5,"Niederösterreich"
"Y15-24","AT13",2013,16.1,"Wien"
"Y15-24","AT2",2013,9.4,"Südösterreich"
"Y15-24","AT21",2013,9.1,"Kärnten"
"Y15-24","AT22",2013,9.6,"Steiermark"
"Y15-24","AT3",2013,6.7,"Westösterreich"
"Y15-24","AT31",2013,7.3,"Oberösterreich"
"Y15-24","AT32",2013,NA,"Salzburg"
"Y15-24","AT33",2013,6.2,"Tirol"
"Y15-24","AT34",2013,NA,"Vorarlberg"
"Y15-24","BE",2013,23.7,"Belgium"
"Y15-24","BE1",2013,39.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2013,39.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2013,16.6,"Vlaams Gewest"
"Y15-24","BE21",2013,19.1,"Prov. Antwerpen"
"Y15-24","BE22",2013,19.8,"Prov. Limburg (BE)"
"Y15-24","BE23",2013,14.4,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2013,16.1,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2013,13.7,"Prov. West-Vlaanderen"
"Y15-24","BE3",2013,32.8,"Région wallonne"
"Y15-24","BE31",2013,29.3,"Prov. Brabant Wallon"
"Y15-24","BE32",2013,40.5,"Prov. Hainaut"
"Y15-24","BE33",2013,26.9,"Prov. Liège"
"Y15-24","BE34",2013,25.9,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2013,32.4,"Prov. Namur"
"Y15-24","BG",2013,28.4,"Bulgaria"
"Y15-24","BG3",2013,31.4,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2013,32,"Severozapaden"
"Y15-24","BG32",2013,29.3,"Severen tsentralen"
"Y15-24","BG33",2013,33,"Severoiztochen"
"Y15-24","BG34",2013,30.7,"Yugoiztochen"
"Y15-24","BG4",2013,25.6,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2013,20.6,"Yugozapaden"
"Y15-24","BG42",2013,34.1,"Yuzhen tsentralen"
"Y15-24","CH",2013,8.5,"Switzerland"
"Y15-24","CH0",2013,8.5,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2013,16,"Région lémanique"
"Y15-24","CH02",2013,7.8,"Espace Mittelland"
"Y15-24","CH03",2013,6.2,"Nordwestschweiz"
"Y15-24","CH04",2013,6.9,"Zürich"
"Y15-24","CH05",2013,6.7,"Ostschweiz"
"Y15-24","CH06",2013,4.3,"Zentralschweiz"
"Y15-24","CH07",2013,16.2,"Ticino"
"Y15-24","CY",2013,38.9,"Cyprus"
"Y15-24","CY0",2013,38.9,"Kypros"
"Y15-24","CY00",2013,38.9,"Kypros"
"Y15-24","CZ",2013,19,"Czech Republic"
"Y15-24","CZ0",2013,19,"Ceská republika"
"Y15-24","CZ01",2013,9.7,"Praha"
"Y15-24","CZ02",2013,14.7,"Strední Cechy"
"Y15-24","CZ03",2013,16.6,"Jihozápad"
"Y15-24","CZ04",2013,24.8,"Severozápad"
"Y15-24","CZ05",2013,19.7,"Severovýchod"
"Y15-24","CZ06",2013,19.4,"Jihovýchod"
"Y15-24","CZ07",2013,21.6,"Strední Morava"
"Y15-24","CZ08",2013,22.4,"Moravskoslezsko"
"Y15-24","DE",2013,7.8,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2013,5.4,"Baden-Württemberg"
"Y15-24","DE11",2013,6,"Stuttgart"
"Y15-24","DE12",2013,5.7,"Karlsruhe"
"Y15-24","DE13",2013,4.7,"Freiburg"
"Y15-24","DE14",2013,4.4,"Tübingen"
"Y15-24","DE2",2013,4.8,"Bayern"
"Y15-24","DE21",2013,4.3,"Oberbayern"
"Y15-24","DE22",2013,NA,"Niederbayern"
"Y15-24","DE23",2013,NA,"Oberpfalz"
"Y15-24","DE24",2013,8,"Oberfranken"
"Y15-24","DE25",2013,4.9,"Mittelfranken"
"Y15-24","DE26",2013,NA,"Unterfranken"
"Y15-24","DE27",2013,4.6,"Schwaben"
"Y15-24","DE3",2013,14.3,"Berlin"
"Y15-24","DE30",2013,14.3,"Berlin"
"Y15-24","DE4",2013,11,"Brandenburg"
"Y15-24","DE40",2013,11,"Brandenburg"
"Y15-24","DE5",2013,NA,"Bremen"
"Y15-24","DE50",2013,NA,"Bremen"
"Y15-24","DE6",2013,7.5,"Hamburg"
"Y15-24","DE60",2013,7.5,"Hamburg"
"Y15-24","DE7",2013,8.1,"Hessen"
"Y15-24","DE71",2013,8.1,"Darmstadt"
"Y15-24","DE72",2013,NA,"Gießen"
"Y15-24","DE73",2013,8.9,"Kassel"
"Y15-24","DE8",2013,11,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2013,11,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2013,7.9,"Niedersachsen"
"Y15-24","DE91",2013,9.5,"Braunschweig"
"Y15-24","DE92",2013,8.6,"Hannover"
"Y15-24","DE93",2013,7.8,"Lüneburg"
"Y15-24","DE94",2013,6.7,"Weser-Ems"
"Y15-24","DEA",2013,9.3,"Nordrhein-Westfalen"
"Y15-24","DEA1",2013,10.1,"Düsseldorf"
"Y15-24","DEA2",2013,8.6,"Köln"
"Y15-24","DEA3",2013,8.5,"Münster"
"Y15-24","DEA4",2013,8.8,"Detmold"
"Y15-24","DEA5",2013,10,"Arnsberg"
"Y15-24","DEB",2013,7.8,"Rheinland-Pfalz"
"Y15-24","DEB1",2013,7,"Koblenz"
"Y15-24","DEB2",2013,NA,"Trier"
"Y15-24","DEB3",2013,9.5,"Rheinhessen-Pfalz"
"Y15-24","DEC",2013,11.9,"Saarland"
"Y15-24","DEC0",2013,11.9,"Saarland"
"Y15-24","DED",2013,10.3,"Sachsen"
"Y15-24","DED2",2013,9.8,"Dresden"
"Y15-24","DED4",2013,9.1,"Chemnitz"
"Y15-24","DED5",2013,12.5,"Leipzig"
"Y15-24","DEE",2013,11.3,"Sachsen-Anhalt"
"Y15-24","DEE0",2013,11.3,"Sachsen-Anhalt"
"Y15-24","DEF",2013,7.1,"Schleswig-Holstein"
"Y15-24","DEF0",2013,7.1,"Schleswig-Holstein"
"Y15-24","DEG",2013,8.7,"Thüringen"
"Y15-24","DEG0",2013,8.7,"Thüringen"
"Y15-24","DK",2013,13.1,"Denmark"
"Y15-24","DK0",2013,13.1,"Danmark"
"Y15-24","DK01",2013,12.7,"Hovedstaden"
"Y15-24","DK02",2013,13.9,"Sjælland"
"Y15-24","DK03",2013,12.8,"Syddanmark"
"Y15-24","DK04",2013,12.7,"Midtjylland"
"Y15-24","DK05",2013,14.4,"Nordjylland"
"Y15-24","EA17",2013,24.4,"Euro area (17 countries)"
"Y15-24","EA18",2013,24.4,"Euro area (18 countries)"
"Y15-24","EA19",2013,24.4,"Euro area (19 countries)"
"Y15-24","EE",2013,18.7,"Estonia"
"Y15-24","EE0",2013,18.7,"Eesti"
"Y15-24","EE00",2013,18.7,"Eesti"
"Y15-24","EL",2013,58.3,"Greece"
"Y15-24","EL3",2013,60.6,"Attiki"
"Y15-24","EL30",2013,60.6,"Attiki"
"Y15-24","EL4",2013,42.9,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2013,46.1,"Voreio Aigaio"
"Y15-24","EL42",2013,37.2,"Notio Aigaio"
"Y15-24","EL43",2013,45.4,"Kriti"
"Y15-24","EL5",2013,62.5,"Voreia Ellada"
"Y15-24","EL51",2013,59.4,"Anatoliki Makedonia, Thraki"
"Y15-24","EL52",2013,62,"Kentriki Makedonia"
"Y15-24","EL53",2013,70.4,"Dytiki Makedonia"
"Y15-24","EL54",2013,67.4,"Ipeiros"
"Y15-24","EL6",2013,58.4,"Kentriki Ellada"
"Y15-24","EL61",2013,57.5,"Thessalia"
"Y15-24","EL62",2013,51.5,"Ionia Nisia"
"Y15-24","EL63",2013,59,"Dytiki Ellada"
"Y15-24","EL64",2013,59.5,"Sterea Ellada"
"Y15-24","EL65",2013,60.3,"Peloponnisos"
"Y15-24","ES",2013,55.5,"Spain"
"Y15-24","ES1",2013,51.3,"Noroeste (ES)"
"Y15-24","ES11",2013,49.9,"Galicia"
"Y15-24","ES12",2013,55,"Principado de Asturias"
"Y15-24","ES13",2013,52.5,"Cantabria"
"Y15-24","ES2",2013,48.2,"Noreste (ES)"
"Y15-24","ES21",2013,46.5,"País Vasco"
"Y15-24","ES22",2013,48.3,"Comunidad Foral de Navarra"
"Y15-24","ES23",2013,48,"La Rioja"
"Y15-24","ES24",2013,50.2,"Aragón"
"Y15-24","ES3",2013,48.8,"Comunidad de Madrid"
"Y15-24","ES30",2013,48.8,"Comunidad de Madrid"
"Y15-24","ES4",2013,57.4,"Centro (ES)"
"Y15-24","ES41",2013,49.7,"Castilla y León"
"Y15-24","ES42",2013,61.5,"Castilla-la Mancha"
"Y15-24","ES43",2013,61.5,"Extremadura"
"Y15-24","ES5",2013,51.9,"Este (ES)"
"Y15-24","ES51",2013,50.2,"Cataluña"
"Y15-24","ES52",2013,56.3,"Comunidad Valenciana"
"Y15-24","ES53",2013,45.2,"Illes Balears"
"Y15-24","ES6",2013,64.1,"Sur (ES)"
"Y15-24","ES61",2013,66,"Andalucía"
"Y15-24","ES62",2013,53.5,"Región de Murcia"
"Y15-24","ES63",2013,73.4,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2013,54,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2013,65.3,"Canarias (ES)"
"Y15-24","ES70",2013,65.3,"Canarias (ES)"
"Y15-24","EU15",2013,23.2,"European Union (15 countries)"
"Y15-24","EU27",2013,23.6,"European Union (27 countries)"
"Y15-24","EU28",2013,23.8,"European Union (28 countries)"
"Y15-24","FI",2013,19.9,"Finland"
"Y15-24","FI1",2013,19.9,"Manner-Suomi"
"Y15-24","FI19",2013,21.9,"Länsi-Suomi"
"Y15-24","FI1B",2013,17.2,"Helsinki-Uusimaa"
"Y15-24","FI1C",2013,20.8,"Etelä-Suomi"
"Y15-24","FI1D",2013,20.8,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2013,NA,"Åland"
"Y15-24","FI20",2013,NA,"Åland"
"Y15-24","FR",2013,25,"France"
"Y15-24","FR1",2013,18.5,"Île de France"
"Y15-24","FR10",2013,18.5,"Île de France"
"Y15-24","FR2",2013,27.6,"Bassin Parisien"
"Y15-24","FR21",2013,30.5,"Champagne-Ardenne"
"Y15-24","FR22",2013,29.3,"Picardie"
"Y15-24","FR23",2013,30.9,"Haute-Normandie"
"Y15-24","FR24",2013,22.1,"Centre (FR)"
"Y15-24","FR25",2013,25.9,"Basse-Normandie"
"Y15-24","FR26",2013,30.4,"Bourgogne"
"Y15-24","FR3",2013,34.9,"Nord - Pas-de-Calais"
"Y15-24","FR30",2013,34.9,"Nord - Pas-de-Calais"
"Y15-24","FR4",2013,26.9,"Est (FR)"
"Y15-24","FR41",2013,27.4,"Lorraine"
"Y15-24","FR42",2013,28.4,"Alsace"
"Y15-24","FR43",2013,22.6,"Franche-Comté"
"Y15-24","FR5",2013,21.7,"Ouest (FR)"
"Y15-24","FR51",2013,20.8,"Pays de la Loire"
"Y15-24","FR52",2013,19.3,"Bretagne"
"Y15-24","FR53",2013,26.5,"Poitou-Charentes"
"Y15-24","FR6",2013,20.7,"Sud-Ouest (FR)"
"Y15-24","FR61",2013,21.9,"Aquitaine"
"Y15-24","FR62",2013,20.5,"Midi-Pyrénées"
"Y15-24","FR63",2013,16.5,"Limousin"
"Y15-24","FR7",2013,20.4,"Centre-Est (FR)"
"Y15-24","FR71",2013,19.5,"Rhône-Alpes"
"Y15-24","FR72",2013,24.8,"Auvergne"
"Y15-24","FR8",2013,28.6,"Méditerranée"
"Y15-24","FR81",2013,36.4,"Languedoc-Roussillon"
"Y15-24","FR82",2013,24.8,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2013,NA,"Corse"
"Y15-24","FRA",2013,57,"Départements d'outre-mer"
"Y15-24","FRA1",2013,58.4,"Guadeloupe"
"Y15-24","FRA2",2013,63.9,"Martinique"
"Y15-24","FRA3",2013,41.1,"Guyane"
"Y15-24","FRA4",2013,57.3,"La Réunion"
"Y15-24","HR",2013,50,"Croatia"
"Y15-24","HR0",2013,50,"Hrvatska"
"Y15-24","HR03",2013,45.2,"Jadranska Hrvatska"
"Y15-24","HR04",2013,51.8,"Kontinentalna Hrvatska"
"Y15-24","HU",2013,26.6,"Hungary"
"Y15-24","HU1",2013,25.2,"Közép-Magyarország"
"Y15-24","HU10",2013,25.2,"Közép-Magyarország"
"Y15-24","HU2",2013,21.6,"Dunántúl"
"Y15-24","HU21",2013,22.7,"Közép-Dunántúl"
"Y15-24","HU22",2013,20.8,"Nyugat-Dunántúl"
"Y15-24","HU23",2013,21.3,"Dél-Dunántúl"
"Y15-24","HU3",2013,31.1,"Alföld és Észak"
"Y15-24","HU31",2013,28.9,"Észak-Magyarország"
"Y15-24","HU32",2013,35.8,"Észak-Alföld"
"Y15-24","HU33",2013,27.3,"Dél-Alföld"
"Y15-24","IE",2013,26.8,"Ireland"
"Y15-24","IE0",2013,26.8,"Éire/Ireland"
"Y15-24","IE01",2013,30.3,"Border, Midland and Western"
"Y15-24","IE02",2013,25.6,"Southern and Eastern"
"Y15-24","IS",2013,10.6,"Iceland"
"Y15-24","IS0",2013,10.6,"Ísland"
"Y15-24","IS00",2013,10.6,"Ísland"
"Y15-24","IT",2013,40,"Italy"
"Y15-24","ITC",2013,34.3,"Nord-Ovest"
"Y15-24","ITC1",2013,40.6,"Piemonte"
"Y15-24","ITC2",2013,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2013,41.2,"Liguria"
"Y15-24","ITC4",2013,30.8,"Lombardia"
"Y15-24","ITF",2013,50.4,"Sud"
"Y15-24","ITF1",2013,36.3,"Abruzzo"
"Y15-24","ITF2",2013,48.6,"Molise"
"Y15-24","ITF3",2013,51.7,"Campania"
"Y15-24","ITF4",2013,49.7,"Puglia"
"Y15-24","ITF5",2013,55.6,"Basilicata"
"Y15-24","ITF6",2013,55.4,"Calabria"
"Y15-24","ITG",2013,54.2,"Isole"
"Y15-24","ITG1",2013,54.3,"Sicilia"
"Y15-24","ITG2",2013,53.7,"Sardegna"
"Y15-24","ITH",2013,27.2,"Nord-Est"
"Y15-24","ITH1",2013,12.1,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2013,23.4,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2013,25.7,"Veneto"
"Y15-24","ITH4",2013,24.5,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2013,33.6,"Emilia-Romagna"
"Y15-24","ITI",2013,39.3,"Centro (IT)"
"Y15-24","ITI1",2013,33.1,"Toscana"
"Y15-24","ITI2",2013,37.2,"Umbria"
"Y15-24","ITI3",2013,36.2,"Marche"
"Y15-24","ITI4",2013,45.1,"Lazio"
"Y15-24","LT",2013,21.9,"Lithuania"
"Y15-24","LT0",2013,21.9,"Lietuva"
"Y15-24","LT00",2013,21.9,"Lietuva"
"Y15-24","LU",2013,15.5,"Luxembourg"
"Y15-24","LU0",2013,15.5,"Luxembourg"
"Y15-24","LU00",2013,15.5,"Luxembourg"
"Y15-24","LV",2013,23.2,"Latvia"
"Y15-24","LV0",2013,23.2,"Latvija"
"Y15-24","LV00",2013,23.2,"Latvija"
"Y15-24","MK",2013,51.9,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2013,51.9,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2013,51.9,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2013,13,"Malta"
"Y15-24","MT0",2013,13,"Malta"
"Y15-24","MT00",2013,13,"Malta"
"Y15-24","NL",2013,13.2,"Netherlands"
"Y15-24","NL1",2013,14.4,"Noord-Nederland"
"Y15-24","NL11",2013,13.9,"Groningen"
"Y15-24","NL12",2013,15.8,"Friesland (NL)"
"Y15-24","NL13",2013,13.1,"Drenthe"
"Y15-24","NL2",2013,13.7,"Oost-Nederland"
"Y15-24","NL21",2013,13.5,"Overijssel"
"Y15-24","NL22",2013,12.6,"Gelderland"
"Y15-24","NL23",2013,19.8,"Flevoland"
"Y15-24","NL3",2013,12.9,"West-Nederland"
"Y15-24","NL31",2013,11.7,"Utrecht"
"Y15-24","NL32",2013,14,"Noord-Holland"
"Y15-24","NL33",2013,13.1,"Zuid-Holland"
"Y15-24","NL34",2013,8.4,"Zeeland"
"Y15-24","NL4",2013,12.6,"Zuid-Nederland"
"Y15-24","NL41",2013,11.7,"Noord-Brabant"
"Y15-24","NL42",2013,14.7,"Limburg (NL)"
"Y15-24","NO",2013,9.1,"Norway"
"Y15-24","NO0",2013,9.1,"Norge"
"Y15-24","NO01",2013,10.3,"Oslo og Akershus"
"Y15-24","NO02",2013,9.2,"Hedmark og Oppland"
"Y15-24","NO03",2013,10.1,"Sør-Østlandet"
"Y15-24","NO04",2013,7.5,"Agder og Rogaland"
"Y15-24","NO05",2013,8.8,"Vestlandet"
"Y15-24","NO06",2013,7,"Trøndelag"
"Y15-24","NO07",2013,10,"Nord-Norge"
"Y15-24","PL",2013,27.3,"Poland"
"Y15-24","PL1",2013,21,"Region Centralny"
"Y15-24","PL11",2013,23.8,"Lódzkie"
"Y15-24","PL12",2013,19.3,"Mazowieckie"
"Y15-24","PL2",2013,27.9,"Region Poludniowy"
"Y15-24","PL21",2013,30.9,"Malopolskie"
"Y15-24","PL22",2013,25.6,"Slaskie"
"Y15-24","PL3",2013,34.3,"Region Wschodni"
"Y15-24","PL31",2013,31,"Lubelskie"
"Y15-24","PL32",2013,43.5,"Podkarpackie"
"Y15-24","PL33",2013,32.2,"Swietokrzyskie"
"Y15-24","PL34",2013,25.8,"Podlaskie"
"Y15-24","PL4",2013,25,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2013,21.9,"Wielkopolskie"
"Y15-24","PL42",2013,32.2,"Zachodniopomorskie"
"Y15-24","PL43",2013,27.8,"Lubuskie"
"Y15-24","PL5",2013,27.9,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2013,30.1,"Dolnoslaskie"
"Y15-24","PL52",2013,21.8,"Opolskie"
"Y15-24","PL6",2013,29.2,"Region Pólnocny"
"Y15-24","PL61",2013,32.3,"Kujawsko-Pomorskie"
"Y15-24","PL62",2013,28.8,"Warminsko-Mazurskie"
"Y15-24","PL63",2013,26.5,"Pomorskie"
"Y15-24","PT",2013,38.1,"Portugal"
"Y15-24","PT1",2013,37.6,"Continente"
"Y15-24","PT11",2013,35.4,"Norte"
"Y15-24","PT15",2013,39.6,"Algarve"
"Y15-24","PT16",2013,31.6,"Centro (PT)"
"Y15-24","PT17",2013,45.3,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2013,39.5,"Alentejo"
"Y15-24","PT2",2013,39.6,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2013,39.6,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2013,51.8,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2013,51.8,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2013,23.7,"Romania"
"Y15-24","RO1",2013,23.3,"Macroregiunea unu"
"Y15-24","RO11",2013,16.4,"Nord-Vest"
"Y15-24","RO12",2013,32.1,"Centru"
"Y15-24","RO2",2013,18.6,"Macroregiunea doi"
"Y15-24","RO21",2013,12.1,"Nord-Est"
"Y15-24","RO22",2013,29.4,"Sud-Est"
"Y15-24","RO3",2013,30,"Macroregiunea trei"
"Y15-24","RO31",2013,32.4,"Sud - Muntenia"
"Y15-24","RO32",2013,25.9,"Bucuresti - Ilfov"
"Y15-24","RO4",2013,23.6,"Macroregiunea patru"
"Y15-24","RO41",2013,23.3,"Sud-Vest Oltenia"
"Y15-24","RO42",2013,24,"Vest"
"Y15-24","SE",2013,23.5,"Sweden"
"Y15-24","SE1",2013,21.7,"Östra Sverige"
"Y15-24","SE11",2013,19.8,"Stockholm"
"Y15-24","SE12",2013,24.1,"Östra Mellansverige"
"Y15-24","SE2",2013,24.8,"Södra Sverige"
"Y15-24","SE21",2013,22.2,"Småland med öarna"
"Y15-24","SE22",2013,27.5,"Sydsverige"
"Y15-24","SE23",2013,24.1,"Västsverige"
"Y15-24","SE3",2013,24.4,"Norra Sverige"
"Y15-24","SE31",2013,26.6,"Norra Mellansverige"
"Y15-24","SE32",2013,23.4,"Mellersta Norrland"
"Y15-24","SE33",2013,21.5,"Övre Norrland"
"Y15-24","SI",2013,21.6,"Slovenia"
"Y15-24","SI0",2013,21.6,"Slovenija"
"Y15-24","SI03",2013,26.2,"Vzhodna Slovenija"
"Y15-24","SI04",2013,16.5,"Zahodna Slovenija"
"Y15-24","SK",2013,33.7,"Slovakia"
"Y15-24","SK0",2013,33.7,"Slovensko"
"Y15-24","SK01",2013,19.7,"Bratislavský kraj"
"Y15-24","SK02",2013,29.5,"Západné Slovensko"
"Y15-24","SK03",2013,35.8,"Stredné Slovensko"
"Y15-24","SK04",2013,39.8,"Východné Slovensko"
"Y15-24","TR",2013,16.9,"Turkey"
"Y15-24","TR1",2013,18.3,"Istanbul"
"Y15-24","TR10",2013,18.3,"Istanbul"
"Y15-24","TR2",2013,14.4,"Bati Marmara"
"Y15-24","TR21",2013,13.3,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2013,15.8,"Balikesir, Çanakkale"
"Y15-24","TR3",2013,18.4,"Ege"
"Y15-24","TR31",2013,25.2,"Izmir"
"Y15-24","TR32",2013,12.8,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2013,12.9,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2013,16.6,"Dogu Marmara"
"Y15-24","TR41",2013,13.2,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2013,20,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2013,16.2,"Bati Anadolu"
"Y15-24","TR51",2013,20.7,"Ankara"
"Y15-24","TR52",2013,7.7,"Konya, Karaman"
"Y15-24","TR6",2013,17.6,"Akdeniz"
"Y15-24","TR61",2013,15,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2013,19.6,"Adana, Mersin"
"Y15-24","TR63",2013,17.3,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2013,14.9,"Orta Anadolu"
"Y15-24","TR71",2013,12.8,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2013,16.1,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2013,14.6,"Bati Karadeniz"
"Y15-24","TR81",2013,15.8,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2013,13.6,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2013,14.4,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2013,20.3,"Dogu Karadeniz"
"Y15-24","TR90",2013,20.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2013,10,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2013,11.2,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2013,9.3,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2013,14,"Ortadogu Anadolu"
"Y15-24","TRB1",2013,11.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2013,16,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2013,18.9,"Güneydogu Anadolu"
"Y15-24","TRC1",2013,10.2,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2013,19.6,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2013,27.6,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2013,20.7,"United Kingdom"
"Y15-24","UKC",2013,26.4,"North East (UK)"
"Y15-24","UKC1",2013,30.2,"Tees Valley and Durham"
"Y15-24","UKC2",2013,23.5,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2013,19.4,"North West (UK)"
"Y15-24","UKD1",2013,12.2,"Cumbria"
"Y15-24","UKD3",2013,22,"Greater Manchester"
"Y15-24","UKD4",2013,19.9,"Lancashire"
"Y15-24","UKD6",2013,15,"Cheshire"
"Y15-24","UKD7",2013,18.3,"Merseyside"
"Y15-24","UKE",2013,23.2,"Yorkshire and The Humber"
"Y15-24","UKE1",2013,21,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2013,13.2,"North Yorkshire"
"Y15-24","UKE3",2013,25.8,"South Yorkshire"
"Y15-24","UKE4",2013,25.2,"West Yorkshire"
"Y15-24","UKF",2013,18.3,"East Midlands (UK)"
"Y15-24","UKF1",2013,19.1,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2013,16.7,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2013,19.4,"Lincolnshire"
"Y15-24","UKG",2013,24.7,"West Midlands (UK)"
"Y15-24","UKG1",2013,15.5,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2013,15.3,"Shropshire and Staffordshire"
"Y15-24","UKG3",2013,33.8,"West Midlands"
"Y15-24","UKH",2013,17.7,"East of England"
"Y15-24","UKH1",2013,18,"East Anglia"
"Y15-24","UKH2",2013,15.7,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2013,18.9,"Essex"
"Y15-24","UKI",2013,25.3,"London"
"Y15-24","UKI3",2013,14,"Inner London - West"
"Y15-24","UKI4",2013,27.9,"Inner London - East"
"Y15-24","UKI5",2013,25.8,"Outer London - East and North East"
"Y15-24","UKI6",2013,26.6,"Outer London - South"
"Y15-24","UKI7",2013,25,"Outer London - West and North West"
"Y15-24","UKJ",2013,17.8,"South East (UK)"
"Y15-24","UKJ1",2013,17.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2013,16.4,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2013,16.6,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2013,21.3,"Kent"
"Y15-24","UKK",2013,17.5,"South West (UK)"
"Y15-24","UKK1",2013,17.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2013,14.6,"Dorset and Somerset"
"Y15-24","UKK3",2013,14.2,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2013,21.4,"Devon"
"Y15-24","UKL",2013,21.1,"Wales"
"Y15-24","UKL1",2013,20.4,"West Wales and The Valleys"
"Y15-24","UKL2",2013,22.3,"East Wales"
"Y15-24","UKM",2013,19.1,"Scotland"
"Y15-24","UKM2",2013,23.1,"Eastern Scotland"
"Y15-24","UKM3",2013,19.2,"South Western Scotland"
"Y15-24","UKM5",2013,NA,"North Eastern Scotland"
"Y15-24","UKM6",2013,14.6,"Highlands and Islands"
"Y15-24","UKN",2013,22.3,"Northern Ireland (UK)"
"Y15-24","UKN0",2013,22.3,"Northern Ireland (UK)"
"Y20-64","AT",2013,5.1,"Austria"
"Y20-64","AT1",2013,6.7,"Ostösterreich"
"Y20-64","AT11",2013,4.1,"Burgenland (AT)"
"Y20-64","AT12",2013,4.5,"Niederösterreich"
"Y20-64","AT13",2013,9,"Wien"
"Y20-64","AT2",2013,4.7,"Südösterreich"
"Y20-64","AT21",2013,5.3,"Kärnten"
"Y20-64","AT22",2013,4.5,"Steiermark"
"Y20-64","AT3",2013,3.5,"Westösterreich"
"Y20-64","AT31",2013,4.2,"Oberösterreich"
"Y20-64","AT32",2013,3,"Salzburg"
"Y20-64","AT33",2013,2.9,"Tirol"
"Y20-64","AT34",2013,3.3,"Vorarlberg"
"Y20-64","BE",2013,8.3,"Belgium"
"Y20-64","BE1",2013,19,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2013,19,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2013,4.9,"Vlaams Gewest"
"Y20-64","BE21",2013,6.1,"Prov. Antwerpen"
"Y20-64","BE22",2013,5.1,"Prov. Limburg (BE)"
"Y20-64","BE23",2013,3.9,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2013,5.4,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2013,3.7,"Prov. West-Vlaanderen"
"Y20-64","BE3",2013,11.1,"Région wallonne"
"Y20-64","BE31",2013,8,"Prov. Brabant Wallon"
"Y20-64","BE32",2013,12.9,"Prov. Hainaut"
"Y20-64","BE33",2013,11.5,"Prov. Liège"
"Y20-64","BE34",2013,7.7,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2013,10.3,"Prov. Namur"
"Y20-64","BG",2013,12.7,"Bulgaria"
"Y20-64","BG3",2013,14.6,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2013,13.7,"Severozapaden"
"Y20-64","BG32",2013,15.2,"Severen tsentralen"
"Y20-64","BG33",2013,16.5,"Severoiztochen"
"Y20-64","BG34",2013,12.9,"Yugoiztochen"
"Y20-64","BG4",2013,11.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2013,9.7,"Yugozapaden"
"Y20-64","BG42",2013,13.2,"Yuzhen tsentralen"
"Y20-64","CH",2013,4.3,"Switzerland"
"Y20-64","CH0",2013,4.3,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2013,6.1,"Région lémanique"
"Y20-64","CH02",2013,3.7,"Espace Mittelland"
"Y20-64","CH03",2013,4.1,"Nordwestschweiz"
"Y20-64","CH04",2013,4.2,"Zürich"
"Y20-64","CH05",2013,3.4,"Ostschweiz"
"Y20-64","CH06",2013,2.7,"Zentralschweiz"
"Y20-64","CH07",2013,6.5,"Ticino"
"Y20-64","CY",2013,15.8,"Cyprus"
"Y20-64","CY0",2013,15.8,"Kypros"
"Y20-64","CY00",2013,15.8,"Kypros"
"Y20-64","CZ",2013,6.8,"Czech Republic"
"Y20-64","CZ0",2013,6.8,"Ceská republika"
"Y20-64","CZ01",2013,3.1,"Praha"
"Y20-64","CZ02",2013,5.1,"Strední Cechy"
"Y20-64","CZ03",2013,5.1,"Jihozápad"
"Y20-64","CZ04",2013,9.5,"Severozápad"
"Y20-64","CZ05",2013,8.1,"Severovýchod"
"Y20-64","CZ06",2013,6.7,"Jihovýchod"
"Y20-64","CZ07",2013,7.9,"Strední Morava"
"Y20-64","CZ08",2013,9.8,"Moravskoslezsko"
"Y20-64","DE",2013,5.2,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2013,3.3,"Baden-Württemberg"
"Y20-64","DE11",2013,3.6,"Stuttgart"
"Y20-64","DE12",2013,3.6,"Karlsruhe"
"Y20-64","DE13",2013,2.8,"Freiburg"
"Y20-64","DE14",2013,2.9,"Tübingen"
"Y20-64","DE2",2013,3,"Bayern"
"Y20-64","DE21",2013,2.5,"Oberbayern"
"Y20-64","DE22",2013,3.3,"Niederbayern"
"Y20-64","DE23",2013,3.4,"Oberpfalz"
"Y20-64","DE24",2013,3.8,"Oberfranken"
"Y20-64","DE25",2013,3.1,"Mittelfranken"
"Y20-64","DE26",2013,3.3,"Unterfranken"
"Y20-64","DE27",2013,3.3,"Schwaben"
"Y20-64","DE3",2013,10.3,"Berlin"
"Y20-64","DE30",2013,10.3,"Berlin"
"Y20-64","DE4",2013,7.3,"Brandenburg"
"Y20-64","DE40",2013,7.3,"Brandenburg"
"Y20-64","DE5",2013,6.9,"Bremen"
"Y20-64","DE50",2013,6.9,"Bremen"
"Y20-64","DE6",2013,4.7,"Hamburg"
"Y20-64","DE60",2013,4.7,"Hamburg"
"Y20-64","DE7",2013,4.3,"Hessen"
"Y20-64","DE71",2013,4.3,"Darmstadt"
"Y20-64","DE72",2013,4.4,"Gießen"
"Y20-64","DE73",2013,4.1,"Kassel"
"Y20-64","DE8",2013,10.1,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2013,10.1,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2013,4.8,"Niedersachsen"
"Y20-64","DE91",2013,6.1,"Braunschweig"
"Y20-64","DE92",2013,5.4,"Hannover"
"Y20-64","DE93",2013,4.2,"Lüneburg"
"Y20-64","DE94",2013,4,"Weser-Ems"
"Y20-64","DEA",2013,5.9,"Nordrhein-Westfalen"
"Y20-64","DEA1",2013,6.3,"Düsseldorf"
"Y20-64","DEA2",2013,5.8,"Köln"
"Y20-64","DEA3",2013,5.2,"Münster"
"Y20-64","DEA4",2013,4.9,"Detmold"
"Y20-64","DEA5",2013,6.5,"Arnsberg"
"Y20-64","DEB",2013,3.9,"Rheinland-Pfalz"
"Y20-64","DEB1",2013,3.6,"Koblenz"
"Y20-64","DEB2",2013,3,"Trier"
"Y20-64","DEB3",2013,4.3,"Rheinhessen-Pfalz"
"Y20-64","DEC",2013,5.9,"Saarland"
"Y20-64","DEC0",2013,5.9,"Saarland"
"Y20-64","DED",2013,7.9,"Sachsen"
"Y20-64","DED2",2013,7.3,"Dresden"
"Y20-64","DED4",2013,7.6,"Chemnitz"
"Y20-64","DED5",2013,9.2,"Leipzig"
"Y20-64","DEE",2013,9.2,"Sachsen-Anhalt"
"Y20-64","DEE0",2013,9.2,"Sachsen-Anhalt"
"Y20-64","DEF",2013,4.9,"Schleswig-Holstein"
"Y20-64","DEF0",2013,4.9,"Schleswig-Holstein"
"Y20-64","DEG",2013,6.1,"Thüringen"
"Y20-64","DEG0",2013,6.1,"Thüringen"
"Y20-64","DK",2013,6.6,"Denmark"
"Y20-64","DK0",2013,6.6,"Danmark"
"Y20-64","DK01",2013,7,"Hovedstaden"
"Y20-64","DK02",2013,6.2,"Sjælland"
"Y20-64","DK03",2013,6.9,"Syddanmark"
"Y20-64","DK04",2013,6,"Midtjylland"
"Y20-64","DK05",2013,5.9,"Nordjylland"
"Y20-64","EA17",2013,11.8,"Euro area (17 countries)"
"Y20-64","EA18",2013,11.8,"Euro area (18 countries)"
"Y20-64","EA19",2013,11.8,"Euro area (19 countries)"
"Y20-64","EE",2013,8.6,"Estonia"
"Y20-64","EE0",2013,8.6,"Eesti"
"Y20-64","EE00",2013,8.6,"Eesti"
"Y20-64","EL",2013,27.3,"Greece"
"Y20-64","EL3",2013,28.3,"Attiki"
"Y20-64","EL30",2013,28.3,"Attiki"
"Y20-64","EL4",2013,23.3,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2013,21.5,"Voreio Aigaio"
"Y20-64","EL42",2013,21.2,"Notio Aigaio"
"Y20-64","EL43",2013,25,"Kriti"
"Y20-64","EL5",2013,29.2,"Voreia Ellada"
"Y20-64","EL51",2013,26.5,"Anatoliki Makedonia, Thraki"
"Y20-64","EL52",2013,30,"Kentriki Makedonia"
"Y20-64","EL53",2013,31.5,"Dytiki Makedonia"
"Y20-64","EL54",2013,27.5,"Ipeiros"
"Y20-64","EL6",2013,25.3,"Kentriki Ellada"
"Y20-64","EL61",2013,25.5,"Thessalia"
"Y20-64","EL62",2013,17.9,"Ionia Nisia"
"Y20-64","EL63",2013,28.1,"Dytiki Ellada"
"Y20-64","EL64",2013,27.9,"Sterea Ellada"
"Y20-64","EL65",2013,22.1,"Peloponnisos"
"Y20-64","ES",2013,25.6,"Spain"
"Y20-64","ES1",2013,22.2,"Noroeste (ES)"
"Y20-64","ES11",2013,22,"Galicia"
"Y20-64","ES12",2013,24,"Principado de Asturias"
"Y20-64","ES13",2013,20.4,"Cantabria"
"Y20-64","ES2",2013,18.1,"Noreste (ES)"
"Y20-64","ES21",2013,16.3,"País Vasco"
"Y20-64","ES22",2013,17.6,"Comunidad Foral de Navarra"
"Y20-64","ES23",2013,19.7,"La Rioja"
"Y20-64","ES24",2013,20.7,"Aragón"
"Y20-64","ES3",2013,19.3,"Comunidad de Madrid"
"Y20-64","ES30",2013,19.3,"Comunidad de Madrid"
"Y20-64","ES4",2013,26.7,"Centro (ES)"
"Y20-64","ES41",2013,21.4,"Castilla y León"
"Y20-64","ES42",2013,29.4,"Castilla-la Mancha"
"Y20-64","ES43",2013,33.4,"Extremadura"
"Y20-64","ES5",2013,24.2,"Este (ES)"
"Y20-64","ES51",2013,22.5,"Cataluña"
"Y20-64","ES52",2013,27.6,"Comunidad Valenciana"
"Y20-64","ES53",2013,21.9,"Illes Balears"
"Y20-64","ES6",2013,34.6,"Sur (ES)"
"Y20-64","ES61",2013,35.7,"Andalucía"
"Y20-64","ES62",2013,28.6,"Región de Murcia"
"Y20-64","ES63",2013,34.2,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2013,32.3,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2013,33.3,"Canarias (ES)"
"Y20-64","ES70",2013,33.3,"Canarias (ES)"
"Y20-64","EU15",2013,10.8,"European Union (15 countries)"
"Y20-64","EU27",2013,10.6,"European Union (27 countries)"
"Y20-64","EU28",2013,10.6,"European Union (28 countries)"
"Y20-64","FI",2013,7.5,"Finland"
"Y20-64","FI1",2013,7.5,"Manner-Suomi"
"Y20-64","FI19",2013,7.9,"Länsi-Suomi"
"Y20-64","FI1B",2013,6,"Helsinki-Uusimaa"
"Y20-64","FI1C",2013,7.8,"Etelä-Suomi"
"Y20-64","FI1D",2013,9,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2013,NA,"Åland"
"Y20-64","FI20",2013,NA,"Åland"
"Y20-64","FR",2013,10,"France"
"Y20-64","FR1",2013,8.9,"Île de France"
"Y20-64","FR10",2013,8.9,"Île de France"
"Y20-64","FR2",2013,10.2,"Bassin Parisien"
"Y20-64","FR21",2013,9.7,"Champagne-Ardenne"
"Y20-64","FR22",2013,10.9,"Picardie"
"Y20-64","FR23",2013,11,"Haute-Normandie"
"Y20-64","FR24",2013,10.2,"Centre (FR)"
"Y20-64","FR25",2013,8.5,"Basse-Normandie"
"Y20-64","FR26",2013,10.2,"Bourgogne"
"Y20-64","FR3",2013,14,"Nord - Pas-de-Calais"
"Y20-64","FR30",2013,14,"Nord - Pas-de-Calais"
"Y20-64","FR4",2013,10.3,"Est (FR)"
"Y20-64","FR41",2013,11.6,"Lorraine"
"Y20-64","FR42",2013,9.1,"Alsace"
"Y20-64","FR43",2013,9.6,"Franche-Comté"
"Y20-64","FR5",2013,8.3,"Ouest (FR)"
"Y20-64","FR51",2013,8.4,"Pays de la Loire"
"Y20-64","FR52",2013,7.6,"Bretagne"
"Y20-64","FR53",2013,9.2,"Poitou-Charentes"
"Y20-64","FR6",2013,8.3,"Sud-Ouest (FR)"
"Y20-64","FR61",2013,8.6,"Aquitaine"
"Y20-64","FR62",2013,8.3,"Midi-Pyrénées"
"Y20-64","FR63",2013,6.7,"Limousin"
"Y20-64","FR7",2013,8.1,"Centre-Est (FR)"
"Y20-64","FR71",2013,8,"Rhône-Alpes"
"Y20-64","FR72",2013,8.5,"Auvergne"
"Y20-64","FR8",2013,11.2,"Méditerranée"
"Y20-64","FR81",2013,12.3,"Languedoc-Roussillon"
"Y20-64","FR82",2013,10.6,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2013,12,"Corse"
"Y20-64","FRA",2013,25.6,"Départements d'outre-mer"
"Y20-64","FRA1",2013,25.9,"Guadeloupe"
"Y20-64","FRA2",2013,22.3,"Martinique"
"Y20-64","FRA3",2013,21.2,"Guyane"
"Y20-64","FRA4",2013,28.1,"La Réunion"
"Y20-64","HR",2013,16.6,"Croatia"
"Y20-64","HR0",2013,16.6,"Hrvatska"
"Y20-64","HR03",2013,14.3,"Jadranska Hrvatska"
"Y20-64","HR04",2013,17.7,"Kontinentalna Hrvatska"
"Y20-64","HU",2013,10,"Hungary"
"Y20-64","HU1",2013,8.6,"Közép-Magyarország"
"Y20-64","HU10",2013,8.6,"Közép-Magyarország"
"Y20-64","HU2",2013,8.3,"Dunántúl"
"Y20-64","HU21",2013,8.6,"Közép-Dunántúl"
"Y20-64","HU22",2013,7.5,"Nyugat-Dunántúl"
"Y20-64","HU23",2013,9,"Dél-Dunántúl"
"Y20-64","HU3",2013,12.5,"Alföld és Észak"
"Y20-64","HU31",2013,12.4,"Észak-Magyarország"
"Y20-64","HU32",2013,14,"Észak-Alföld"
"Y20-64","HU33",2013,10.8,"Dél-Alföld"
"Y20-64","IE",2013,12.9,"Ireland"
"Y20-64","IE0",2013,12.9,"Éire/Ireland"
"Y20-64","IE01",2013,14.1,"Border, Midland and Western"
"Y20-64","IE02",2013,12.4,"Southern and Eastern"
"Y20-64","IS",2013,4.8,"Iceland"
"Y20-64","IS0",2013,4.8,"Ísland"
"Y20-64","IS00",2013,4.8,"Ísland"
"Y20-64","IT",2013,11.9,"Italy"
"Y20-64","ITC",2013,8.6,"Nord-Ovest"
"Y20-64","ITC1",2013,10.2,"Piemonte"
"Y20-64","ITC2",2013,8.1,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2013,9.8,"Liguria"
"Y20-64","ITC4",2013,7.8,"Lombardia"
"Y20-64","ITF",2013,19.2,"Sud"
"Y20-64","ITF1",2013,11.2,"Abruzzo"
"Y20-64","ITF2",2013,15.4,"Molise"
"Y20-64","ITF3",2013,21,"Campania"
"Y20-64","ITF4",2013,19.3,"Puglia"
"Y20-64","ITF5",2013,15,"Basilicata"
"Y20-64","ITF6",2013,22,"Calabria"
"Y20-64","ITG",2013,19.6,"Isole"
"Y20-64","ITG1",2013,20.6,"Sicilia"
"Y20-64","ITG2",2013,17.1,"Sardegna"
"Y20-64","ITH",2013,7.5,"Nord-Est"
"Y20-64","ITH1",2013,4.2,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2013,6.3,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2013,7.4,"Veneto"
"Y20-64","ITH4",2013,7.6,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2013,8.1,"Emilia-Romagna"
"Y20-64","ITI",2013,10.5,"Centro (IT)"
"Y20-64","ITI1",2013,8.5,"Toscana"
"Y20-64","ITI2",2013,10.1,"Umbria"
"Y20-64","ITI3",2013,10.8,"Marche"
"Y20-64","ITI4",2013,11.7,"Lazio"
"Y20-64","LT",2013,11.9,"Lithuania"
"Y20-64","LT0",2013,11.9,"Lietuva"
"Y20-64","LT00",2013,11.9,"Lietuva"
"Y20-64","LU",2013,5.7,"Luxembourg"
"Y20-64","LU0",2013,5.7,"Luxembourg"
"Y20-64","LU00",2013,5.7,"Luxembourg"
"Y20-64","LV",2013,11.9,"Latvia"
"Y20-64","LV0",2013,11.9,"Latvija"
"Y20-64","LV00",2013,11.9,"Latvija"
"Y20-64","MK",2013,28.5,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2013,28.5,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2013,28.5,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2013,5.7,"Malta"
"Y20-64","MT0",2013,5.7,"Malta"
"Y20-64","MT00",2013,5.7,"Malta"
"Y20-64","NL",2013,6.7,"Netherlands"
"Y20-64","NL1",2013,7.3,"Noord-Nederland"
"Y20-64","NL11",2013,7.6,"Groningen"
"Y20-64","NL12",2013,7.7,"Friesland (NL)"
"Y20-64","NL13",2013,6.4,"Drenthe"
"Y20-64","NL2",2013,6.6,"Oost-Nederland"
"Y20-64","NL21",2013,6.7,"Overijssel"
"Y20-64","NL22",2013,6,"Gelderland"
"Y20-64","NL23",2013,9.1,"Flevoland"
"Y20-64","NL3",2013,6.8,"West-Nederland"
"Y20-64","NL31",2013,5.8,"Utrecht"
"Y20-64","NL32",2013,6.5,"Noord-Holland"
"Y20-64","NL33",2013,7.5,"Zuid-Holland"
"Y20-64","NL34",2013,4.3,"Zeeland"
"Y20-64","NL4",2013,6.3,"Zuid-Nederland"
"Y20-64","NL41",2013,6,"Noord-Brabant"
"Y20-64","NL42",2013,6.8,"Limburg (NL)"
"Y20-64","NO",2013,3,"Norway"
"Y20-64","NO0",2013,3,"Norge"
"Y20-64","NO01",2013,3.5,"Oslo og Akershus"
"Y20-64","NO02",2013,2.8,"Hedmark og Oppland"
"Y20-64","NO03",2013,3.4,"Sør-Østlandet"
"Y20-64","NO04",2013,2.9,"Agder og Rogaland"
"Y20-64","NO05",2013,2.7,"Vestlandet"
"Y20-64","NO06",2013,2.5,"Trøndelag"
"Y20-64","NO07",2013,2.7,"Nord-Norge"
"Y20-64","PL",2013,10.2,"Poland"
"Y20-64","PL1",2013,9.1,"Region Centralny"
"Y20-64","PL11",2013,11.1,"Lódzkie"
"Y20-64","PL12",2013,7.9,"Mazowieckie"
"Y20-64","PL2",2013,10.1,"Region Poludniowy"
"Y20-64","PL21",2013,10.8,"Malopolskie"
"Y20-64","PL22",2013,9.6,"Slaskie"
"Y20-64","PL3",2013,12,"Region Wschodni"
"Y20-64","PL31",2013,10.3,"Lubelskie"
"Y20-64","PL32",2013,14.5,"Podkarpackie"
"Y20-64","PL33",2013,13,"Swietokrzyskie"
"Y20-64","PL34",2013,9.9,"Podlaskie"
"Y20-64","PL4",2013,9.1,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2013,8.6,"Wielkopolskie"
"Y20-64","PL42",2013,9.9,"Zachodniopomorskie"
"Y20-64","PL43",2013,9.5,"Lubuskie"
"Y20-64","PL5",2013,10.7,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2013,11.1,"Dolnoslaskie"
"Y20-64","PL52",2013,9.4,"Opolskie"
"Y20-64","PL6",2013,11,"Region Pólnocny"
"Y20-64","PL61",2013,12.2,"Kujawsko-Pomorskie"
"Y20-64","PL62",2013,11.1,"Warminsko-Mazurskie"
"Y20-64","PL63",2013,9.9,"Pomorskie"
"Y20-64","PT",2013,16.5,"Portugal"
"Y20-64","PT1",2013,16.5,"Continente"
"Y20-64","PT11",2013,17.4,"Norte"
"Y20-64","PT15",2013,17,"Algarve"
"Y20-64","PT16",2013,12.1,"Centro (PT)"
"Y20-64","PT17",2013,18.5,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2013,17.2,"Alentejo"
"Y20-64","PT2",2013,16.8,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2013,16.8,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2013,18.2,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2013,18.2,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2013,7.1,"Romania"
"Y20-64","RO1",2013,6.3,"Macroregiunea unu"
"Y20-64","RO11",2013,4,"Nord-Vest"
"Y20-64","RO12",2013,9.1,"Centru"
"Y20-64","RO2",2013,6.5,"Macroregiunea doi"
"Y20-64","RO21",2013,4.6,"Nord-Est"
"Y20-64","RO22",2013,9.3,"Sud-Est"
"Y20-64","RO3",2013,8.8,"Macroregiunea trei"
"Y20-64","RO31",2013,9.5,"Sud - Muntenia"
"Y20-64","RO32",2013,8,"Bucuresti - Ilfov"
"Y20-64","RO4",2013,6.2,"Macroregiunea patru"
"Y20-64","RO41",2013,7.3,"Sud-Vest Oltenia"
"Y20-64","RO42",2013,4.9,"Vest"
"Y20-64","SE",2013,7.1,"Sweden"
"Y20-64","SE1",2013,6.7,"Östra Sverige"
"Y20-64","SE11",2013,5.9,"Stockholm"
"Y20-64","SE12",2013,7.9,"Östra Mellansverige"
"Y20-64","SE2",2013,7.5,"Södra Sverige"
"Y20-64","SE21",2013,6.2,"Småland med öarna"
"Y20-64","SE22",2013,8.9,"Sydsverige"
"Y20-64","SE23",2013,7.1,"Västsverige"
"Y20-64","SE3",2013,7.2,"Norra Sverige"
"Y20-64","SE31",2013,8.1,"Norra Mellansverige"
"Y20-64","SE32",2013,6.1,"Mellersta Norrland"
"Y20-64","SE33",2013,6.5,"Övre Norrland"
"Y20-64","SI",2013,10.2,"Slovenia"
"Y20-64","SI0",2013,10.2,"Slovenija"
"Y20-64","SI03",2013,11.5,"Vzhodna Slovenija"
"Y20-64","SI04",2013,8.8,"Zahodna Slovenija"
"Y20-64","SK",2013,13.9,"Slovakia"
"Y20-64","SK0",2013,13.9,"Slovensko"
"Y20-64","SK01",2013,6.3,"Bratislavský kraj"
"Y20-64","SK02",2013,11.5,"Západné Slovensko"
"Y20-64","SK03",2013,16.3,"Stredné Slovensko"
"Y20-64","SK04",2013,18,"Východné Slovensko"
"Y20-64","TR",2013,8.6,"Turkey"
"Y20-64","TR1",2013,10.2,"Istanbul"
"Y20-64","TR10",2013,10.2,"Istanbul"
"Y20-64","TR2",2013,5.9,"Bati Marmara"
"Y20-64","TR21",2013,6.3,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2013,5.5,"Balikesir, Çanakkale"
"Y20-64","TR3",2013,9.1,"Ege"
"Y20-64","TR31",2013,13.9,"Izmir"
"Y20-64","TR32",2013,6,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2013,5.2,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2013,7.4,"Dogu Marmara"
"Y20-64","TR41",2013,5.9,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2013,8.9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2013,7.3,"Bati Anadolu"
"Y20-64","TR51",2013,8.7,"Ankara"
"Y20-64","TR52",2013,3.8,"Konya, Karaman"
"Y20-64","TR6",2013,9.7,"Akdeniz"
"Y20-64","TR61",2013,7,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2013,11.2,"Adana, Mersin"
"Y20-64","TR63",2013,11.2,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2013,7.3,"Orta Anadolu"
"Y20-64","TR71",2013,5.5,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2013,8.4,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2013,5.7,"Bati Karadeniz"
"Y20-64","TR81",2013,6.2,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2013,5.5,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2013,5.6,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2013,6,"Dogu Karadeniz"
"Y20-64","TR90",2013,6,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2013,5.8,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2013,6.1,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2013,5.5,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2013,7.1,"Ortadogu Anadolu"
"Y20-64","TRB1",2013,5.7,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2013,8.7,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2013,12.7,"Güneydogu Anadolu"
"Y20-64","TRC1",2013,6,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2013,15.9,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2013,18.2,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2013,6.7,"United Kingdom"
"Y20-64","UKC",2013,8.8,"North East (UK)"
"Y20-64","UKC1",2013,9.1,"Tees Valley and Durham"
"Y20-64","UKC2",2013,8.6,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2013,7.2,"North West (UK)"
"Y20-64","UKD1",2013,4.6,"Cumbria"
"Y20-64","UKD3",2013,8.5,"Greater Manchester"
"Y20-64","UKD4",2013,6.3,"Lancashire"
"Y20-64","UKD6",2013,4.4,"Cheshire"
"Y20-64","UKD7",2013,8.1,"Merseyside"
"Y20-64","UKE",2013,7.5,"Yorkshire and The Humber"
"Y20-64","UKE1",2013,7.6,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2013,4,"North Yorkshire"
"Y20-64","UKE3",2013,8.7,"South Yorkshire"
"Y20-64","UKE4",2013,8,"West Yorkshire"
"Y20-64","UKF",2013,6.7,"East Midlands (UK)"
"Y20-64","UKF1",2013,6.6,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2013,7.3,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2013,5.7,"Lincolnshire"
"Y20-64","UKG",2013,8.3,"West Midlands (UK)"
"Y20-64","UKG1",2013,4.6,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2013,5.5,"Shropshire and Staffordshire"
"Y20-64","UKG3",2013,11.8,"West Midlands"
"Y20-64","UKH",2013,5.3,"East of England"
"Y20-64","UKH1",2013,5.5,"East Anglia"
"Y20-64","UKH2",2013,4.9,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2013,5.6,"Essex"
"Y20-64","UKI",2013,7.8,"London"
"Y20-64","UKI3",2013,6.5,"Inner London - West"
"Y20-64","UKI4",2013,8.9,"Inner London - East"
"Y20-64","UKI5",2013,8.3,"Outer London - East and North East"
"Y20-64","UKI6",2013,6.3,"Outer London - South"
"Y20-64","UKI7",2013,7.6,"Outer London - West and North West"
"Y20-64","UKJ",2013,5,"South East (UK)"
"Y20-64","UKJ1",2013,4.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2013,4.6,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2013,4.9,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2013,6.5,"Kent"
"Y20-64","UKK",2013,5.4,"South West (UK)"
"Y20-64","UKK1",2013,5.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2013,4.8,"Dorset and Somerset"
"Y20-64","UKK3",2013,5.5,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2013,6.2,"Devon"
"Y20-64","UKL",2013,6.9,"Wales"
"Y20-64","UKL1",2013,7.2,"West Wales and The Valleys"
"Y20-64","UKL2",2013,6.5,"East Wales"
"Y20-64","UKM",2013,6.2,"Scotland"
"Y20-64","UKM2",2013,6.1,"Eastern Scotland"
"Y20-64","UKM3",2013,7.2,"South Western Scotland"
"Y20-64","UKM5",2013,4.3,"North Eastern Scotland"
"Y20-64","UKM6",2013,5,"Highlands and Islands"
"Y20-64","UKN",2013,7.2,"Northern Ireland (UK)"
"Y20-64","UKN0",2013,7.2,"Northern Ireland (UK)"
"Y_GE15","AT",2013,5.3,"Austria"
"Y_GE15","AT1",2013,7,"Ostösterreich"
"Y_GE15","AT11",2013,4.3,"Burgenland (AT)"
"Y_GE15","AT12",2013,5,"Niederösterreich"
"Y_GE15","AT13",2013,9.2,"Wien"
"Y_GE15","AT2",2013,4.9,"Südösterreich"
"Y_GE15","AT21",2013,5.5,"Kärnten"
"Y_GE15","AT22",2013,4.7,"Steiermark"
"Y_GE15","AT3",2013,3.7,"Westösterreich"
"Y_GE15","AT31",2013,4.3,"Oberösterreich"
"Y_GE15","AT32",2013,3.2,"Salzburg"
"Y_GE15","AT33",2013,3.1,"Tirol"
"Y_GE15","AT34",2013,3.6,"Vorarlberg"
"Y_GE15","BE",2013,8.4,"Belgium"
"Y_GE15","BE1",2013,19.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2013,19.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2013,5,"Vlaams Gewest"
"Y_GE15","BE21",2013,6.2,"Prov. Antwerpen"
"Y_GE15","BE22",2013,5.5,"Prov. Limburg (BE)"
"Y_GE15","BE23",2013,4,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2013,5.5,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2013,3.9,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2013,11.3,"Région wallonne"
"Y_GE15","BE31",2013,8.2,"Prov. Brabant Wallon"
"Y_GE15","BE32",2013,13.2,"Prov. Hainaut"
"Y_GE15","BE33",2013,11.7,"Prov. Liège"
"Y_GE15","BE34",2013,7.9,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2013,10.4,"Prov. Namur"
"Y_GE15","BG",2013,12.9,"Bulgaria"
"Y_GE15","BG3",2013,14.8,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2013,14,"Severozapaden"
"Y_GE15","BG32",2013,15.3,"Severen tsentralen"
"Y_GE15","BG33",2013,16.8,"Severoiztochen"
"Y_GE15","BG34",2013,13,"Yugoiztochen"
"Y_GE15","BG4",2013,11.2,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2013,9.8,"Yugozapaden"
"Y_GE15","BG42",2013,13.5,"Yuzhen tsentralen"
"Y_GE15","CH",2013,4.4,"Switzerland"
"Y_GE15","CH0",2013,4.4,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2013,6.6,"Région lémanique"
"Y_GE15","CH02",2013,3.8,"Espace Mittelland"
"Y_GE15","CH03",2013,4.1,"Nordwestschweiz"
"Y_GE15","CH04",2013,4.2,"Zürich"
"Y_GE15","CH05",2013,3.6,"Ostschweiz"
"Y_GE15","CH06",2013,2.6,"Zentralschweiz"
"Y_GE15","CH07",2013,6.8,"Ticino"
"Y_GE15","CY",2013,15.9,"Cyprus"
"Y_GE15","CY0",2013,15.9,"Kypros"
"Y_GE15","CY00",2013,15.9,"Kypros"
"Y_GE15","CZ",2013,7,"Czech Republic"
"Y_GE15","CZ0",2013,7,"Ceská republika"
"Y_GE15","CZ01",2013,3.1,"Praha"
"Y_GE15","CZ02",2013,5.2,"Strední Cechy"
"Y_GE15","CZ03",2013,5.2,"Jihozápad"
"Y_GE15","CZ04",2013,9.6,"Severozápad"
"Y_GE15","CZ05",2013,8.3,"Severovýchod"
"Y_GE15","CZ06",2013,6.8,"Jihovýchod"
"Y_GE15","CZ07",2013,8,"Strední Morava"
"Y_GE15","CZ08",2013,9.9,"Moravskoslezsko"
"Y_GE15","DE",2013,5.2,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2013,3.3,"Baden-Württemberg"
"Y_GE15","DE11",2013,3.6,"Stuttgart"
"Y_GE15","DE12",2013,3.6,"Karlsruhe"
"Y_GE15","DE13",2013,2.9,"Freiburg"
"Y_GE15","DE14",2013,2.9,"Tübingen"
"Y_GE15","DE2",2013,3,"Bayern"
"Y_GE15","DE21",2013,2.5,"Oberbayern"
"Y_GE15","DE22",2013,3.2,"Niederbayern"
"Y_GE15","DE23",2013,3.4,"Oberpfalz"
"Y_GE15","DE24",2013,3.9,"Oberfranken"
"Y_GE15","DE25",2013,3.1,"Mittelfranken"
"Y_GE15","DE26",2013,3.3,"Unterfranken"
"Y_GE15","DE27",2013,3.3,"Schwaben"
"Y_GE15","DE3",2013,10.4,"Berlin"
"Y_GE15","DE30",2013,10.4,"Berlin"
"Y_GE15","DE4",2013,7.3,"Brandenburg"
"Y_GE15","DE40",2013,7.3,"Brandenburg"
"Y_GE15","DE5",2013,7,"Bremen"
"Y_GE15","DE50",2013,7,"Bremen"
"Y_GE15","DE6",2013,4.7,"Hamburg"
"Y_GE15","DE60",2013,4.7,"Hamburg"
"Y_GE15","DE7",2013,4.3,"Hessen"
"Y_GE15","DE71",2013,4.3,"Darmstadt"
"Y_GE15","DE72",2013,4.5,"Gießen"
"Y_GE15","DE73",2013,4.3,"Kassel"
"Y_GE15","DE8",2013,10,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2013,10,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2013,4.9,"Niedersachsen"
"Y_GE15","DE91",2013,6.2,"Braunschweig"
"Y_GE15","DE92",2013,5.4,"Hannover"
"Y_GE15","DE93",2013,4.3,"Lüneburg"
"Y_GE15","DE94",2013,4,"Weser-Ems"
"Y_GE15","DEA",2013,5.9,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2013,6.3,"Düsseldorf"
"Y_GE15","DEA2",2013,5.8,"Köln"
"Y_GE15","DEA3",2013,5.1,"Münster"
"Y_GE15","DEA4",2013,5,"Detmold"
"Y_GE15","DEA5",2013,6.5,"Arnsberg"
"Y_GE15","DEB",2013,4,"Rheinland-Pfalz"
"Y_GE15","DEB1",2013,3.8,"Koblenz"
"Y_GE15","DEB2",2013,3,"Trier"
"Y_GE15","DEB3",2013,4.4,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2013,5.9,"Saarland"
"Y_GE15","DEC0",2013,5.9,"Saarland"
"Y_GE15","DED",2013,7.8,"Sachsen"
"Y_GE15","DED2",2013,7.2,"Dresden"
"Y_GE15","DED4",2013,7.4,"Chemnitz"
"Y_GE15","DED5",2013,9.2,"Leipzig"
"Y_GE15","DEE",2013,9.1,"Sachsen-Anhalt"
"Y_GE15","DEE0",2013,9.1,"Sachsen-Anhalt"
"Y_GE15","DEF",2013,4.9,"Schleswig-Holstein"
"Y_GE15","DEF0",2013,4.9,"Schleswig-Holstein"
"Y_GE15","DEG",2013,6,"Thüringen"
"Y_GE15","DEG0",2013,6,"Thüringen"
"Y_GE15","DK",2013,7,"Denmark"
"Y_GE15","DK0",2013,7,"Danmark"
"Y_GE15","DK01",2013,7.4,"Hovedstaden"
"Y_GE15","DK02",2013,6.8,"Sjælland"
"Y_GE15","DK03",2013,7.2,"Syddanmark"
"Y_GE15","DK04",2013,6.5,"Midtjylland"
"Y_GE15","DK05",2013,6.4,"Nordjylland"
"Y_GE15","EA17",2013,12,"Euro area (17 countries)"
"Y_GE15","EA18",2013,12,"Euro area (18 countries)"
"Y_GE15","EA19",2013,12,"Euro area (19 countries)"
"Y_GE15","EE",2013,8.6,"Estonia"
"Y_GE15","EE0",2013,8.6,"Eesti"
"Y_GE15","EE00",2013,8.6,"Eesti"
"Y_GE15","EL",2013,27.5,"Greece"
"Y_GE15","EL3",2013,28.7,"Attiki"
"Y_GE15","EL30",2013,28.7,"Attiki"
"Y_GE15","EL4",2013,23.4,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2013,22,"Voreio Aigaio"
"Y_GE15","EL42",2013,21.3,"Notio Aigaio"
"Y_GE15","EL43",2013,24.9,"Kriti"
"Y_GE15","EL5",2013,29.3,"Voreia Ellada"
"Y_GE15","EL51",2013,26.8,"Anatoliki Makedonia, Thraki"
"Y_GE15","EL52",2013,30.2,"Kentriki Makedonia"
"Y_GE15","EL53",2013,31.6,"Dytiki Makedonia"
"Y_GE15","EL54",2013,27.4,"Ipeiros"
"Y_GE15","EL6",2013,25.4,"Kentriki Ellada"
"Y_GE15","EL61",2013,25.4,"Thessalia"
"Y_GE15","EL62",2013,18.1,"Ionia Nisia"
"Y_GE15","EL63",2013,28.4,"Dytiki Ellada"
"Y_GE15","EL64",2013,28.2,"Sterea Ellada"
"Y_GE15","EL65",2013,21.9,"Peloponnisos"
"Y_GE15","ES",2013,26.1,"Spain"
"Y_GE15","ES1",2013,22.3,"Noroeste (ES)"
"Y_GE15","ES11",2013,22,"Galicia"
"Y_GE15","ES12",2013,24.1,"Principado de Asturias"
"Y_GE15","ES13",2013,20.4,"Cantabria"
"Y_GE15","ES2",2013,18.5,"Noreste (ES)"
"Y_GE15","ES21",2013,16.6,"País Vasco"
"Y_GE15","ES22",2013,17.9,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2013,20,"La Rioja"
"Y_GE15","ES24",2013,21.4,"Aragón"
"Y_GE15","ES3",2013,19.8,"Comunidad de Madrid"
"Y_GE15","ES30",2013,19.8,"Comunidad de Madrid"
"Y_GE15","ES4",2013,27.1,"Centro (ES)"
"Y_GE15","ES41",2013,21.7,"Castilla y León"
"Y_GE15","ES42",2013,30,"Castilla-la Mancha"
"Y_GE15","ES43",2013,33.9,"Extremadura"
"Y_GE15","ES5",2013,24.8,"Este (ES)"
"Y_GE15","ES51",2013,23.1,"Cataluña"
"Y_GE15","ES52",2013,28,"Comunidad Valenciana"
"Y_GE15","ES53",2013,22.3,"Illes Balears"
"Y_GE15","ES6",2013,35.1,"Sur (ES)"
"Y_GE15","ES61",2013,36.2,"Andalucía"
"Y_GE15","ES62",2013,29,"Región de Murcia"
"Y_GE15","ES63",2013,34.8,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2013,32.5,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2013,33.7,"Canarias (ES)"
"Y_GE15","ES70",2013,33.7,"Canarias (ES)"
"Y_GE15","EU15",2013,11.1,"European Union (15 countries)"
"Y_GE15","EU27",2013,10.8,"European Union (27 countries)"
"Y_GE15","EU28",2013,10.9,"European Union (28 countries)"
"Y_GE15","FI",2013,8.2,"Finland"
"Y_GE15","FI1",2013,8.2,"Manner-Suomi"
"Y_GE15","FI19",2013,8.5,"Länsi-Suomi"
"Y_GE15","FI1B",2013,6.7,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2013,8.4,"Etelä-Suomi"
"Y_GE15","FI1D",2013,9.9,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2013,NA,"Åland"
"Y_GE15","FI20",2013,NA,"Åland"
"Y_GE15","FR",2013,10.3,"France"
"Y_GE15","FR1",2013,9,"Île de France"
"Y_GE15","FR10",2013,9,"Île de France"
"Y_GE15","FR2",2013,10.7,"Bassin Parisien"
"Y_GE15","FR21",2013,10.5,"Champagne-Ardenne"
"Y_GE15","FR22",2013,11.5,"Picardie"
"Y_GE15","FR23",2013,11.5,"Haute-Normandie"
"Y_GE15","FR24",2013,10.5,"Centre (FR)"
"Y_GE15","FR25",2013,9.1,"Basse-Normandie"
"Y_GE15","FR26",2013,10.6,"Bourgogne"
"Y_GE15","FR3",2013,14.7,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2013,14.7,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2013,10.7,"Est (FR)"
"Y_GE15","FR41",2013,12.1,"Lorraine"
"Y_GE15","FR42",2013,9.7,"Alsace"
"Y_GE15","FR43",2013,9.5,"Franche-Comté"
"Y_GE15","FR5",2013,8.7,"Ouest (FR)"
"Y_GE15","FR51",2013,8.8,"Pays de la Loire"
"Y_GE15","FR52",2013,8,"Bretagne"
"Y_GE15","FR53",2013,9.9,"Poitou-Charentes"
"Y_GE15","FR6",2013,8.6,"Sud-Ouest (FR)"
"Y_GE15","FR61",2013,8.9,"Aquitaine"
"Y_GE15","FR62",2013,8.6,"Midi-Pyrénées"
"Y_GE15","FR63",2013,6.9,"Limousin"
"Y_GE15","FR7",2013,8.5,"Centre-Est (FR)"
"Y_GE15","FR71",2013,8.4,"Rhône-Alpes"
"Y_GE15","FR72",2013,8.9,"Auvergne"
"Y_GE15","FR8",2013,11.5,"Méditerranée"
"Y_GE15","FR81",2013,12.9,"Languedoc-Roussillon"
"Y_GE15","FR82",2013,10.8,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2013,12.3,"Corse"
"Y_GE15","FRA",2013,26.2,"Départements d'outre-mer"
"Y_GE15","FRA1",2013,26.2,"Guadeloupe"
"Y_GE15","FRA2",2013,22.8,"Martinique"
"Y_GE15","FRA3",2013,21.3,"Guyane"
"Y_GE15","FRA4",2013,28.9,"La Réunion"
"Y_GE15","HR",2013,17.3,"Croatia"
"Y_GE15","HR0",2013,17.3,"Hrvatska"
"Y_GE15","HR03",2013,15,"Jadranska Hrvatska"
"Y_GE15","HR04",2013,18.3,"Kontinentalna Hrvatska"
"Y_GE15","HU",2013,10.2,"Hungary"
"Y_GE15","HU1",2013,8.7,"Közép-Magyarország"
"Y_GE15","HU10",2013,8.7,"Közép-Magyarország"
"Y_GE15","HU2",2013,8.5,"Dunántúl"
"Y_GE15","HU21",2013,8.7,"Közép-Dunántúl"
"Y_GE15","HU22",2013,7.7,"Nyugat-Dunántúl"
"Y_GE15","HU23",2013,9.3,"Dél-Dunántúl"
"Y_GE15","HU3",2013,12.7,"Alföld és Észak"
"Y_GE15","HU31",2013,12.6,"Észak-Magyarország"
"Y_GE15","HU32",2013,14.2,"Észak-Alföld"
"Y_GE15","HU33",2013,11,"Dél-Alföld"
"Y_GE15","IE",2013,13,"Ireland"
"Y_GE15","IE0",2013,13,"Éire/Ireland"
"Y_GE15","IE01",2013,14.2,"Border, Midland and Western"
"Y_GE15","IE02",2013,12.6,"Southern and Eastern"
"Y_GE15","IS",2013,5.4,"Iceland"
"Y_GE15","IS0",2013,5.4,"Ísland"
"Y_GE15","IS00",2013,5.4,"Ísland"
"Y_GE15","IT",2013,12.1,"Italy"
"Y_GE15","ITC",2013,8.9,"Nord-Ovest"
"Y_GE15","ITC1",2013,10.5,"Piemonte"
"Y_GE15","ITC2",2013,8.3,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2013,9.8,"Liguria"
"Y_GE15","ITC4",2013,8,"Lombardia"
"Y_GE15","ITF",2013,19.5,"Sud"
"Y_GE15","ITF1",2013,11.3,"Abruzzo"
"Y_GE15","ITF2",2013,15.6,"Molise"
"Y_GE15","ITF3",2013,21.5,"Campania"
"Y_GE15","ITF4",2013,19.7,"Puglia"
"Y_GE15","ITF5",2013,15.2,"Basilicata"
"Y_GE15","ITF6",2013,22.3,"Calabria"
"Y_GE15","ITG",2013,20,"Isole"
"Y_GE15","ITG1",2013,21,"Sicilia"
"Y_GE15","ITG2",2013,17.5,"Sardegna"
"Y_GE15","ITH",2013,7.7,"Nord-Est"
"Y_GE15","ITH1",2013,4.4,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2013,6.5,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2013,7.6,"Veneto"
"Y_GE15","ITH4",2013,7.7,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2013,8.4,"Emilia-Romagna"
"Y_GE15","ITI",2013,10.7,"Centro (IT)"
"Y_GE15","ITI1",2013,8.7,"Toscana"
"Y_GE15","ITI2",2013,10.3,"Umbria"
"Y_GE15","ITI3",2013,10.9,"Marche"
"Y_GE15","ITI4",2013,12,"Lazio"
"Y_GE15","LT",2013,11.8,"Lithuania"
"Y_GE15","LT0",2013,11.8,"Lietuva"
"Y_GE15","LT00",2013,11.8,"Lietuva"
"Y_GE15","LU",2013,5.8,"Luxembourg"
"Y_GE15","LU0",2013,5.8,"Luxembourg"
"Y_GE15","LU00",2013,5.8,"Luxembourg"
"Y_GE15","LV",2013,11.9,"Latvia"
"Y_GE15","LV0",2013,11.9,"Latvija"
"Y_GE15","LV00",2013,11.9,"Latvija"
"Y_GE15","MK",2013,29,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2013,29,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2013,29,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2013,6.4,"Malta"
"Y_GE15","MT0",2013,6.4,"Malta"
"Y_GE15","MT00",2013,6.4,"Malta"
"Y_GE15","NL",2013,7.2,"Netherlands"
"Y_GE15","NL1",2013,8,"Noord-Nederland"
"Y_GE15","NL11",2013,8.2,"Groningen"
"Y_GE15","NL12",2013,8.3,"Friesland (NL)"
"Y_GE15","NL13",2013,7.1,"Drenthe"
"Y_GE15","NL2",2013,7.2,"Oost-Nederland"
"Y_GE15","NL21",2013,7.2,"Overijssel"
"Y_GE15","NL22",2013,6.6,"Gelderland"
"Y_GE15","NL23",2013,9.9,"Flevoland"
"Y_GE15","NL3",2013,7.3,"West-Nederland"
"Y_GE15","NL31",2013,6.4,"Utrecht"
"Y_GE15","NL32",2013,7.2,"Noord-Holland"
"Y_GE15","NL33",2013,7.9,"Zuid-Holland"
"Y_GE15","NL34",2013,5,"Zeeland"
"Y_GE15","NL4",2013,6.9,"Zuid-Nederland"
"Y_GE15","NL41",2013,6.7,"Noord-Brabant"
"Y_GE15","NL42",2013,7.4,"Limburg (NL)"
"Y_GE15","NO",2013,3.4,"Norway"
"Y_GE15","NO0",2013,3.4,"Norge"
"Y_GE15","NO01",2013,3.9,"Oslo og Akershus"
"Y_GE15","NO02",2013,2.9,"Hedmark og Oppland"
"Y_GE15","NO03",2013,3.9,"Sør-Østlandet"
"Y_GE15","NO04",2013,3.2,"Agder og Rogaland"
"Y_GE15","NO05",2013,3.1,"Vestlandet"
"Y_GE15","NO06",2013,2.6,"Trøndelag"
"Y_GE15","NO07",2013,3.2,"Nord-Norge"
"Y_GE15","PL",2013,10.3,"Poland"
"Y_GE15","PL1",2013,9.1,"Region Centralny"
"Y_GE15","PL11",2013,11.1,"Lódzkie"
"Y_GE15","PL12",2013,8,"Mazowieckie"
"Y_GE15","PL2",2013,10.2,"Region Poludniowy"
"Y_GE15","PL21",2013,10.9,"Malopolskie"
"Y_GE15","PL22",2013,9.7,"Slaskie"
"Y_GE15","PL3",2013,12,"Region Wschodni"
"Y_GE15","PL31",2013,10.3,"Lubelskie"
"Y_GE15","PL32",2013,14.4,"Podkarpackie"
"Y_GE15","PL33",2013,13,"Swietokrzyskie"
"Y_GE15","PL34",2013,9.9,"Podlaskie"
"Y_GE15","PL4",2013,9.3,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2013,8.8,"Wielkopolskie"
"Y_GE15","PL42",2013,10.1,"Zachodniopomorskie"
"Y_GE15","PL43",2013,9.7,"Lubuskie"
"Y_GE15","PL5",2013,10.8,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2013,11.3,"Dolnoslaskie"
"Y_GE15","PL52",2013,9.4,"Opolskie"
"Y_GE15","PL6",2013,11.2,"Region Pólnocny"
"Y_GE15","PL61",2013,12.4,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2013,11.4,"Warminsko-Mazurskie"
"Y_GE15","PL63",2013,10,"Pomorskie"
"Y_GE15","PT",2013,16.2,"Portugal"
"Y_GE15","PT1",2013,16.1,"Continente"
"Y_GE15","PT11",2013,17.1,"Norte"
"Y_GE15","PT15",2013,16.9,"Algarve"
"Y_GE15","PT16",2013,11.4,"Centro (PT)"
"Y_GE15","PT17",2013,18.5,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2013,16.9,"Alentejo"
"Y_GE15","PT2",2013,17,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2013,17,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2013,18.1,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2013,18.1,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2013,7.1,"Romania"
"Y_GE15","RO1",2013,6.5,"Macroregiunea unu"
"Y_GE15","RO11",2013,4.1,"Nord-Vest"
"Y_GE15","RO12",2013,9.5,"Centru"
"Y_GE15","RO2",2013,6.5,"Macroregiunea doi"
"Y_GE15","RO21",2013,4.4,"Nord-Est"
"Y_GE15","RO22",2013,9.5,"Sud-Est"
"Y_GE15","RO3",2013,8.9,"Macroregiunea trei"
"Y_GE15","RO31",2013,9.5,"Sud - Muntenia"
"Y_GE15","RO32",2013,8,"Bucuresti - Ilfov"
"Y_GE15","RO4",2013,6.2,"Macroregiunea patru"
"Y_GE15","RO41",2013,7,"Sud-Vest Oltenia"
"Y_GE15","RO42",2013,5.2,"Vest"
"Y_GE15","SE",2013,8.1,"Sweden"
"Y_GE15","SE1",2013,7.7,"Östra Sverige"
"Y_GE15","SE11",2013,6.9,"Stockholm"
"Y_GE15","SE12",2013,8.8,"Östra Mellansverige"
"Y_GE15","SE2",2013,8.5,"Södra Sverige"
"Y_GE15","SE21",2013,7.1,"Småland med öarna"
"Y_GE15","SE22",2013,9.9,"Sydsverige"
"Y_GE15","SE23",2013,8,"Västsverige"
"Y_GE15","SE3",2013,8,"Norra Sverige"
"Y_GE15","SE31",2013,8.8,"Norra Mellansverige"
"Y_GE15","SE32",2013,7.2,"Mellersta Norrland"
"Y_GE15","SE33",2013,7.2,"Övre Norrland"
"Y_GE15","SI",2013,10.1,"Slovenia"
"Y_GE15","SI0",2013,10.1,"Slovenija"
"Y_GE15","SI03",2013,11.3,"Vzhodna Slovenija"
"Y_GE15","SI04",2013,8.7,"Zahodna Slovenija"
"Y_GE15","SK",2013,14.2,"Slovakia"
"Y_GE15","SK0",2013,14.2,"Slovensko"
"Y_GE15","SK01",2013,6.4,"Bratislavský kraj"
"Y_GE15","SK02",2013,11.7,"Západné Slovensko"
"Y_GE15","SK03",2013,16.8,"Stredné Slovensko"
"Y_GE15","SK04",2013,18.5,"Východné Slovensko"
"Y_GE15","TR",2013,8.7,"Turkey"
"Y_GE15","TR1",2013,10.6,"Istanbul"
"Y_GE15","TR10",2013,10.6,"Istanbul"
"Y_GE15","TR2",2013,6,"Bati Marmara"
"Y_GE15","TR21",2013,6.4,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2013,5.6,"Balikesir, Çanakkale"
"Y_GE15","TR3",2013,9.3,"Ege"
"Y_GE15","TR31",2013,14.3,"Izmir"
"Y_GE15","TR32",2013,6,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2013,5.2,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2013,7.5,"Dogu Marmara"
"Y_GE15","TR41",2013,6,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2013,9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2013,7.5,"Bati Anadolu"
"Y_GE15","TR51",2013,9,"Ankara"
"Y_GE15","TR52",2013,3.8,"Konya, Karaman"
"Y_GE15","TR6",2013,9.8,"Akdeniz"
"Y_GE15","TR61",2013,7.2,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2013,11.3,"Adana, Mersin"
"Y_GE15","TR63",2013,10.8,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2013,7.3,"Orta Anadolu"
"Y_GE15","TR71",2013,5.5,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2013,8.4,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2013,5.7,"Bati Karadeniz"
"Y_GE15","TR81",2013,6.2,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2013,5.6,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2013,5.5,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2013,6,"Dogu Karadeniz"
"Y_GE15","TR90",2013,6,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2013,5.9,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2013,6.1,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2013,5.6,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2013,7.3,"Ortadogu Anadolu"
"Y_GE15","TRB1",2013,5.7,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2013,9.2,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2013,13.1,"Güneydogu Anadolu"
"Y_GE15","TRC1",2013,6.2,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2013,16,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2013,19.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2013,7.5,"United Kingdom"
"Y_GE15","UKC",2013,10,"North East (UK)"
"Y_GE15","UKC1",2013,10.9,"Tees Valley and Durham"
"Y_GE15","UKC2",2013,9.2,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2013,8,"North West (UK)"
"Y_GE15","UKD1",2013,5.1,"Cumbria"
"Y_GE15","UKD3",2013,9.4,"Greater Manchester"
"Y_GE15","UKD4",2013,7.2,"Lancashire"
"Y_GE15","UKD6",2013,5.2,"Cheshire"
"Y_GE15","UKD7",2013,8.9,"Merseyside"
"Y_GE15","UKE",2013,8.7,"Yorkshire and The Humber"
"Y_GE15","UKE1",2013,8.3,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2013,4.4,"North Yorkshire"
"Y_GE15","UKE3",2013,10.5,"South Yorkshire"
"Y_GE15","UKE4",2013,9.3,"West Yorkshire"
"Y_GE15","UKF",2013,7.3,"East Midlands (UK)"
"Y_GE15","UKF1",2013,7.2,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2013,7.8,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2013,6.4,"Lincolnshire"
"Y_GE15","UKG",2013,9.1,"West Midlands (UK)"
"Y_GE15","UKG1",2013,5.1,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2013,6.2,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2013,13,"West Midlands"
"Y_GE15","UKH",2013,6,"East of England"
"Y_GE15","UKH1",2013,6.2,"East Anglia"
"Y_GE15","UKH2",2013,5.6,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2013,6.3,"Essex"
"Y_GE15","UKI",2013,8.6,"London"
"Y_GE15","UKI3",2013,6.8,"Inner London - West"
"Y_GE15","UKI4",2013,9.8,"Inner London - East"
"Y_GE15","UKI5",2013,9.5,"Outer London - East and North East"
"Y_GE15","UKI6",2013,7.4,"Outer London - South"
"Y_GE15","UKI7",2013,8.4,"Outer London - West and North West"
"Y_GE15","UKJ",2013,5.8,"South East (UK)"
"Y_GE15","UKJ1",2013,5.2,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2013,5.5,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2013,5.7,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2013,7.6,"Kent"
"Y_GE15","UKK",2013,6.1,"South West (UK)"
"Y_GE15","UKK1",2013,6.2,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2013,5.4,"Dorset and Somerset"
"Y_GE15","UKK3",2013,5.6,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2013,7,"Devon"
"Y_GE15","UKL",2013,7.6,"Wales"
"Y_GE15","UKL1",2013,7.8,"West Wales and The Valleys"
"Y_GE15","UKL2",2013,7.4,"East Wales"
"Y_GE15","UKM",2013,7.2,"Scotland"
"Y_GE15","UKM2",2013,7.3,"Eastern Scotland"
"Y_GE15","UKM3",2013,8.2,"South Western Scotland"
"Y_GE15","UKM5",2013,4.8,"North Eastern Scotland"
"Y_GE15","UKM6",2013,5.6,"Highlands and Islands"
"Y_GE15","UKN",2013,7.5,"Northern Ireland (UK)"
"Y_GE15","UKN0",2013,7.5,"Northern Ireland (UK)"
"Y_GE25","AT",2013,4.7,"Austria"
"Y_GE25","AT1",2013,6.1,"Ostösterreich"
"Y_GE25","AT11",2013,3.7,"Burgenland (AT)"
"Y_GE25","AT12",2013,4.1,"Niederösterreich"
"Y_GE25","AT13",2013,8.3,"Wien"
"Y_GE25","AT2",2013,4.2,"Südösterreich"
"Y_GE25","AT21",2013,4.9,"Kärnten"
"Y_GE25","AT22",2013,3.9,"Steiermark"
"Y_GE25","AT3",2013,3.2,"Westösterreich"
"Y_GE25","AT31",2013,3.8,"Oberösterreich"
"Y_GE25","AT32",2013,2.9,"Salzburg"
"Y_GE25","AT33",2013,2.6,"Tirol"
"Y_GE25","AT34",2013,3,"Vorarlberg"
"Y_GE25","BE",2013,7,"Belgium"
"Y_GE25","BE1",2013,17.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2013,17.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2013,4,"Vlaams Gewest"
"Y_GE25","BE21",2013,5,"Prov. Antwerpen"
"Y_GE25","BE22",2013,4.1,"Prov. Limburg (BE)"
"Y_GE25","BE23",2013,3,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2013,4.7,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2013,2.9,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2013,9.3,"Région wallonne"
"Y_GE25","BE31",2013,6.7,"Prov. Brabant Wallon"
"Y_GE25","BE32",2013,10.6,"Prov. Hainaut"
"Y_GE25","BE33",2013,10.2,"Prov. Liège"
"Y_GE25","BE34",2013,5.9,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2013,8.3,"Prov. Namur"
"Y_GE25","BG",2013,11.8,"Bulgaria"
"Y_GE25","BG3",2013,13.6,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2013,12.8,"Severozapaden"
"Y_GE25","BG32",2013,14.4,"Severen tsentralen"
"Y_GE25","BG33",2013,15.4,"Severoiztochen"
"Y_GE25","BG34",2013,11.9,"Yugoiztochen"
"Y_GE25","BG4",2013,10.2,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2013,9,"Yugozapaden"
"Y_GE25","BG42",2013,12,"Yuzhen tsentralen"
"Y_GE25","CH",2013,3.7,"Switzerland"
"Y_GE25","CH0",2013,3.7,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2013,5.2,"Région lémanique"
"Y_GE25","CH02",2013,3.2,"Espace Mittelland"
"Y_GE25","CH03",2013,3.8,"Nordwestschweiz"
"Y_GE25","CH04",2013,3.8,"Zürich"
"Y_GE25","CH05",2013,3,"Ostschweiz"
"Y_GE25","CH06",2013,2.4,"Zentralschweiz"
"Y_GE25","CH07",2013,5.7,"Ticino"
"Y_GE25","CY",2013,13.5,"Cyprus"
"Y_GE25","CY0",2013,13.5,"Kypros"
"Y_GE25","CY00",2013,13.5,"Kypros"
"Y_GE25","CZ",2013,6.1,"Czech Republic"
"Y_GE25","CZ0",2013,6.1,"Ceská republika"
"Y_GE25","CZ01",2013,2.8,"Praha"
"Y_GE25","CZ02",2013,4.5,"Strední Cechy"
"Y_GE25","CZ03",2013,4.4,"Jihozápad"
"Y_GE25","CZ04",2013,8.4,"Severozápad"
"Y_GE25","CZ05",2013,7.3,"Severovýchod"
"Y_GE25","CZ06",2013,5.8,"Jihovýchod"
"Y_GE25","CZ07",2013,7.1,"Strední Morava"
"Y_GE25","CZ08",2013,8.9,"Moravskoslezsko"
"Y_GE25","DE",2013,4.9,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2013,3.1,"Baden-Württemberg"
"Y_GE25","DE11",2013,3.3,"Stuttgart"
"Y_GE25","DE12",2013,3.3,"Karlsruhe"
"Y_GE25","DE13",2013,2.7,"Freiburg"
"Y_GE25","DE14",2013,2.7,"Tübingen"
"Y_GE25","DE2",2013,2.8,"Bayern"
"Y_GE25","DE21",2013,2.3,"Oberbayern"
"Y_GE25","DE22",2013,3,"Niederbayern"
"Y_GE25","DE23",2013,3.3,"Oberpfalz"
"Y_GE25","DE24",2013,3.4,"Oberfranken"
"Y_GE25","DE25",2013,2.9,"Mittelfranken"
"Y_GE25","DE26",2013,3,"Unterfranken"
"Y_GE25","DE27",2013,3.1,"Schwaben"
"Y_GE25","DE3",2013,10,"Berlin"
"Y_GE25","DE30",2013,10,"Berlin"
"Y_GE25","DE4",2013,7,"Brandenburg"
"Y_GE25","DE40",2013,7,"Brandenburg"
"Y_GE25","DE5",2013,6.4,"Bremen"
"Y_GE25","DE50",2013,6.4,"Bremen"
"Y_GE25","DE6",2013,4.4,"Hamburg"
"Y_GE25","DE60",2013,4.4,"Hamburg"
"Y_GE25","DE7",2013,3.9,"Hessen"
"Y_GE25","DE71",2013,3.9,"Darmstadt"
"Y_GE25","DE72",2013,4.2,"Gießen"
"Y_GE25","DE73",2013,3.7,"Kassel"
"Y_GE25","DE8",2013,10,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2013,10,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2013,4.5,"Niedersachsen"
"Y_GE25","DE91",2013,5.9,"Braunschweig"
"Y_GE25","DE92",2013,5.1,"Hannover"
"Y_GE25","DE93",2013,3.9,"Lüneburg"
"Y_GE25","DE94",2013,3.6,"Weser-Ems"
"Y_GE25","DEA",2013,5.5,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2013,5.9,"Düsseldorf"
"Y_GE25","DEA2",2013,5.5,"Köln"
"Y_GE25","DEA3",2013,4.6,"Münster"
"Y_GE25","DEA4",2013,4.6,"Detmold"
"Y_GE25","DEA5",2013,6.1,"Arnsberg"
"Y_GE25","DEB",2013,3.5,"Rheinland-Pfalz"
"Y_GE25","DEB1",2013,3.3,"Koblenz"
"Y_GE25","DEB2",2013,2.9,"Trier"
"Y_GE25","DEB3",2013,3.8,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2013,5.3,"Saarland"
"Y_GE25","DEC0",2013,5.3,"Saarland"
"Y_GE25","DED",2013,7.6,"Sachsen"
"Y_GE25","DED2",2013,7,"Dresden"
"Y_GE25","DED4",2013,7.3,"Chemnitz"
"Y_GE25","DED5",2013,8.9,"Leipzig"
"Y_GE25","DEE",2013,8.9,"Sachsen-Anhalt"
"Y_GE25","DEE0",2013,8.9,"Sachsen-Anhalt"
"Y_GE25","DEF",2013,4.6,"Schleswig-Holstein"
"Y_GE25","DEF0",2013,4.6,"Schleswig-Holstein"
"Y_GE25","DEG",2013,5.8,"Thüringen"
"Y_GE25","DEG0",2013,5.8,"Thüringen"
"Y_GE25","DK",2013,5.9,"Denmark"
"Y_GE25","DK0",2013,5.9,"Danmark"
"Y_GE25","DK01",2013,6.5,"Hovedstaden"
"Y_GE25","DK02",2013,5.7,"Sjælland"
"Y_GE25","DK03",2013,6.2,"Syddanmark"
"Y_GE25","DK04",2013,5.3,"Midtjylland"
"Y_GE25","DK05",2013,4.9,"Nordjylland"
"Y_GE25","EA17",2013,10.7,"Euro area (17 countries)"
"Y_GE25","EA18",2013,10.7,"Euro area (18 countries)"
"Y_GE25","EA19",2013,10.7,"Euro area (19 countries)"
"Y_GE25","EE",2013,7.6,"Estonia"
"Y_GE25","EE0",2013,7.6,"Eesti"
"Y_GE25","EE00",2013,7.6,"Eesti"
"Y_GE25","EL",2013,25.3,"Greece"
"Y_GE25","EL3",2013,26.6,"Attiki"
"Y_GE25","EL30",2013,26.6,"Attiki"
"Y_GE25","EL4",2013,21.8,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2013,19.4,"Voreio Aigaio"
"Y_GE25","EL42",2013,19.9,"Notio Aigaio"
"Y_GE25","EL43",2013,23.4,"Kriti"
"Y_GE25","EL5",2013,27.1,"Voreia Ellada"
"Y_GE25","EL51",2013,24.1,"Anatoliki Makedonia, Thraki"
"Y_GE25","EL52",2013,28.1,"Kentriki Makedonia"
"Y_GE25","EL53",2013,29.3,"Dytiki Makedonia"
"Y_GE25","EL54",2013,24.9,"Ipeiros"
"Y_GE25","EL6",2013,22.9,"Kentriki Ellada"
"Y_GE25","EL61",2013,22.9,"Thessalia"
"Y_GE25","EL62",2013,15.8,"Ionia Nisia"
"Y_GE25","EL63",2013,26,"Dytiki Ellada"
"Y_GE25","EL64",2013,25.3,"Sterea Ellada"
"Y_GE25","EL65",2013,19.7,"Peloponnisos"
"Y_GE25","ES",2013,23.7,"Spain"
"Y_GE25","ES1",2013,20.6,"Noroeste (ES)"
"Y_GE25","ES11",2013,20.3,"Galicia"
"Y_GE25","ES12",2013,22.5,"Principado de Asturias"
"Y_GE25","ES13",2013,18.8,"Cantabria"
"Y_GE25","ES2",2013,16.6,"Noreste (ES)"
"Y_GE25","ES21",2013,15,"País Vasco"
"Y_GE25","ES22",2013,16,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2013,18.2,"La Rioja"
"Y_GE25","ES24",2013,19.2,"Aragón"
"Y_GE25","ES3",2013,17.7,"Comunidad de Madrid"
"Y_GE25","ES30",2013,17.7,"Comunidad de Madrid"
"Y_GE25","ES4",2013,24.7,"Centro (ES)"
"Y_GE25","ES41",2013,19.9,"Castilla y León"
"Y_GE25","ES42",2013,27,"Castilla-la Mancha"
"Y_GE25","ES43",2013,31.1,"Extremadura"
"Y_GE25","ES5",2013,22.5,"Este (ES)"
"Y_GE25","ES51",2013,20.8,"Cataluña"
"Y_GE25","ES52",2013,25.7,"Comunidad Valenciana"
"Y_GE25","ES53",2013,20.4,"Illes Balears"
"Y_GE25","ES6",2013,32.4,"Sur (ES)"
"Y_GE25","ES61",2013,33.4,"Andalucía"
"Y_GE25","ES62",2013,26.7,"Región de Murcia"
"Y_GE25","ES63",2013,31.2,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2013,29.9,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2013,31,"Canarias (ES)"
"Y_GE25","ES70",2013,31,"Canarias (ES)"
"Y_GE25","EU15",2013,9.7,"European Union (15 countries)"
"Y_GE25","EU27",2013,9.4,"European Union (27 countries)"
"Y_GE25","EU28",2013,9.5,"European Union (28 countries)"
"Y_GE25","FI",2013,6.5,"Finland"
"Y_GE25","FI1",2013,6.6,"Manner-Suomi"
"Y_GE25","FI19",2013,6.6,"Länsi-Suomi"
"Y_GE25","FI1B",2013,5.3,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2013,6.8,"Etelä-Suomi"
"Y_GE25","FI1D",2013,8.2,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2013,NA,"Åland"
"Y_GE25","FI20",2013,NA,"Åland"
"Y_GE25","FR",2013,8.8,"France"
"Y_GE25","FR1",2013,8.1,"Île de France"
"Y_GE25","FR10",2013,8.1,"Île de France"
"Y_GE25","FR2",2013,8.8,"Bassin Parisien"
"Y_GE25","FR21",2013,8.1,"Champagne-Ardenne"
"Y_GE25","FR22",2013,9.6,"Picardie"
"Y_GE25","FR23",2013,9.3,"Haute-Normandie"
"Y_GE25","FR24",2013,9.2,"Centre (FR)"
"Y_GE25","FR25",2013,7.2,"Basse-Normandie"
"Y_GE25","FR26",2013,8.8,"Bourgogne"
"Y_GE25","FR3",2013,12.1,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2013,12.1,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2013,8.8,"Est (FR)"
"Y_GE25","FR41",2013,10.3,"Lorraine"
"Y_GE25","FR42",2013,7.4,"Alsace"
"Y_GE25","FR43",2013,8.3,"Franche-Comté"
"Y_GE25","FR5",2013,7.2,"Ouest (FR)"
"Y_GE25","FR51",2013,7.3,"Pays de la Loire"
"Y_GE25","FR52",2013,6.9,"Bretagne"
"Y_GE25","FR53",2013,7.7,"Poitou-Charentes"
"Y_GE25","FR6",2013,7.4,"Sud-Ouest (FR)"
"Y_GE25","FR61",2013,7.6,"Aquitaine"
"Y_GE25","FR62",2013,7.5,"Midi-Pyrénées"
"Y_GE25","FR63",2013,5.9,"Limousin"
"Y_GE25","FR7",2013,7.1,"Centre-Est (FR)"
"Y_GE25","FR71",2013,7.1,"Rhône-Alpes"
"Y_GE25","FR72",2013,7.2,"Auvergne"
"Y_GE25","FR8",2013,9.9,"Méditerranée"
"Y_GE25","FR81",2013,10.7,"Languedoc-Roussillon"
"Y_GE25","FR82",2013,9.5,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2013,10.4,"Corse"
"Y_GE25","FRA",2013,22.5,"Départements d'outre-mer"
"Y_GE25","FRA1",2013,23.3,"Guadeloupe"
"Y_GE25","FRA2",2013,19.2,"Martinique"
"Y_GE25","FRA3",2013,18.8,"Guyane"
"Y_GE25","FRA4",2013,24.7,"La Réunion"
"Y_GE25","HR",2013,14.4,"Croatia"
"Y_GE25","HR0",2013,14.4,"Hrvatska"
"Y_GE25","HR03",2013,12.6,"Jadranska Hrvatska"
"Y_GE25","HR04",2013,15.2,"Kontinentalna Hrvatska"
"Y_GE25","HU",2013,8.9,"Hungary"
"Y_GE25","HU1",2013,7.7,"Közép-Magyarország"
"Y_GE25","HU10",2013,7.7,"Közép-Magyarország"
"Y_GE25","HU2",2013,7.5,"Dunántúl"
"Y_GE25","HU21",2013,7.6,"Közép-Dunántúl"
"Y_GE25","HU22",2013,6.5,"Nyugat-Dunántúl"
"Y_GE25","HU23",2013,8.4,"Dél-Dunántúl"
"Y_GE25","HU3",2013,11,"Alföld és Észak"
"Y_GE25","HU31",2013,11.1,"Észak-Magyarország"
"Y_GE25","HU32",2013,12.3,"Észak-Alföld"
"Y_GE25","HU33",2013,9.5,"Dél-Alföld"
"Y_GE25","IE",2013,11.5,"Ireland"
"Y_GE25","IE0",2013,11.5,"Éire/Ireland"
"Y_GE25","IE01",2013,12.4,"Border, Midland and Western"
"Y_GE25","IE02",2013,11.2,"Southern and Eastern"
"Y_GE25","IS",2013,4.3,"Iceland"
"Y_GE25","IS0",2013,4.3,"Ísland"
"Y_GE25","IS00",2013,4.3,"Ísland"
"Y_GE25","IT",2013,10.2,"Italy"
"Y_GE25","ITC",2013,7.3,"Nord-Ovest"
"Y_GE25","ITC1",2013,8.6,"Piemonte"
"Y_GE25","ITC2",2013,6.8,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2013,8.2,"Liguria"
"Y_GE25","ITC4",2013,6.5,"Lombardia"
"Y_GE25","ITF",2013,16.9,"Sud"
"Y_GE25","ITF1",2013,9.7,"Abruzzo"
"Y_GE25","ITF2",2013,13.2,"Molise"
"Y_GE25","ITF3",2013,18.6,"Campania"
"Y_GE25","ITF4",2013,17.1,"Puglia"
"Y_GE25","ITF5",2013,12.7,"Basilicata"
"Y_GE25","ITF6",2013,19.3,"Calabria"
"Y_GE25","ITG",2013,17.1,"Isole"
"Y_GE25","ITG1",2013,18,"Sicilia"
"Y_GE25","ITG2",2013,14.9,"Sardegna"
"Y_GE25","ITH",2013,6.5,"Nord-Est"
"Y_GE25","ITH1",2013,3.6,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2013,5.3,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2013,6.4,"Veneto"
"Y_GE25","ITH4",2013,6.8,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2013,7,"Emilia-Romagna"
"Y_GE25","ITI",2013,9,"Centro (IT)"
"Y_GE25","ITI1",2013,7.2,"Toscana"
"Y_GE25","ITI2",2013,8.6,"Umbria"
"Y_GE25","ITI3",2013,9.4,"Marche"
"Y_GE25","ITI4",2013,10.1,"Lazio"
"Y_GE25","LT",2013,10.8,"Lithuania"
"Y_GE25","LT0",2013,10.8,"Lietuva"
"Y_GE25","LT00",2013,10.8,"Lietuva"
"Y_GE25","LU",2013,5.2,"Luxembourg"
"Y_GE25","LU0",2013,5.2,"Luxembourg"
"Y_GE25","LU00",2013,5.2,"Luxembourg"
"Y_GE25","LV",2013,10.7,"Latvia"
"Y_GE25","LV0",2013,10.7,"Latvija"
"Y_GE25","LV00",2013,10.7,"Latvija"
"Y_GE25","MK",2013,26.3,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2013,26.3,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2013,26.3,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2013,5.2,"Malta"
"Y_GE25","MT0",2013,5.2,"Malta"
"Y_GE25","MT00",2013,5.2,"Malta"
"Y_GE25","NL",2013,6.1,"Netherlands"
"Y_GE25","NL1",2013,6.8,"Noord-Nederland"
"Y_GE25","NL11",2013,7.1,"Groningen"
"Y_GE25","NL12",2013,7,"Friesland (NL)"
"Y_GE25","NL13",2013,6.1,"Drenthe"
"Y_GE25","NL2",2013,5.9,"Oost-Nederland"
"Y_GE25","NL21",2013,6,"Overijssel"
"Y_GE25","NL22",2013,5.4,"Gelderland"
"Y_GE25","NL23",2013,8.1,"Flevoland"
"Y_GE25","NL3",2013,6.2,"West-Nederland"
"Y_GE25","NL31",2013,5.3,"Utrecht"
"Y_GE25","NL32",2013,6,"Noord-Holland"
"Y_GE25","NL33",2013,7,"Zuid-Holland"
"Y_GE25","NL34",2013,4.4,"Zeeland"
"Y_GE25","NL4",2013,5.8,"Zuid-Nederland"
"Y_GE25","NL41",2013,5.7,"Noord-Brabant"
"Y_GE25","NL42",2013,6.1,"Limburg (NL)"
"Y_GE25","NO",2013,2.5,"Norway"
"Y_GE25","NO0",2013,2.5,"Norge"
"Y_GE25","NO01",2013,3.1,"Oslo og Akershus"
"Y_GE25","NO02",2013,2,"Hedmark og Oppland"
"Y_GE25","NO03",2013,2.9,"Sør-Østlandet"
"Y_GE25","NO04",2013,2.4,"Agder og Rogaland"
"Y_GE25","NO05",2013,2.1,"Vestlandet"
"Y_GE25","NO06",2013,1.9,"Trøndelag"
"Y_GE25","NO07",2013,2,"Nord-Norge"
"Y_GE25","PL",2013,8.7,"Poland"
"Y_GE25","PL1",2013,8.1,"Region Centralny"
"Y_GE25","PL11",2013,10,"Lódzkie"
"Y_GE25","PL12",2013,7.1,"Mazowieckie"
"Y_GE25","PL2",2013,8.4,"Region Poludniowy"
"Y_GE25","PL21",2013,8.6,"Malopolskie"
"Y_GE25","PL22",2013,8.2,"Slaskie"
"Y_GE25","PL3",2013,10,"Region Wschodni"
"Y_GE25","PL31",2013,8.5,"Lubelskie"
"Y_GE25","PL32",2013,11.6,"Podkarpackie"
"Y_GE25","PL33",2013,11.2,"Swietokrzyskie"
"Y_GE25","PL34",2013,8.5,"Podlaskie"
"Y_GE25","PL4",2013,7.7,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2013,7.3,"Wielkopolskie"
"Y_GE25","PL42",2013,8.1,"Zachodniopomorskie"
"Y_GE25","PL43",2013,8.2,"Lubuskie"
"Y_GE25","PL5",2013,9.3,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2013,9.7,"Dolnoslaskie"
"Y_GE25","PL52",2013,8.2,"Opolskie"
"Y_GE25","PL6",2013,9.5,"Region Pólnocny"
"Y_GE25","PL61",2013,10.3,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2013,9.9,"Warminsko-Mazurskie"
"Y_GE25","PL63",2013,8.5,"Pomorskie"
"Y_GE25","PT",2013,14.4,"Portugal"
"Y_GE25","PT1",2013,14.4,"Continente"
"Y_GE25","PT11",2013,15.5,"Norte"
"Y_GE25","PT15",2013,15.2,"Algarve"
"Y_GE25","PT16",2013,10,"Centro (PT)"
"Y_GE25","PT17",2013,16.4,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2013,15.2,"Alentejo"
"Y_GE25","PT2",2013,14.3,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2013,14.3,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2013,15.1,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2013,15.1,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2013,5.7,"Romania"
"Y_GE25","RO1",2013,5.1,"Macroregiunea unu"
"Y_GE25","RO11",2013,3,"Nord-Vest"
"Y_GE25","RO12",2013,7.7,"Centru"
"Y_GE25","RO2",2013,5.4,"Macroregiunea doi"
"Y_GE25","RO21",2013,3.7,"Nord-Est"
"Y_GE25","RO22",2013,7.8,"Sud-Est"
"Y_GE25","RO3",2013,7.2,"Macroregiunea trei"
"Y_GE25","RO31",2013,7.4,"Sud - Muntenia"
"Y_GE25","RO32",2013,6.9,"Bucuresti - Ilfov"
"Y_GE25","RO4",2013,4.9,"Macroregiunea patru"
"Y_GE25","RO41",2013,5.8,"Sud-Vest Oltenia"
"Y_GE25","RO42",2013,3.9,"Vest"
"Y_GE25","SE",2013,5.7,"Sweden"
"Y_GE25","SE1",2013,5.6,"Östra Sverige"
"Y_GE25","SE11",2013,5.1,"Stockholm"
"Y_GE25","SE12",2013,6.3,"Östra Mellansverige"
"Y_GE25","SE2",2013,5.9,"Södra Sverige"
"Y_GE25","SE21",2013,4.6,"Småland med öarna"
"Y_GE25","SE22",2013,7.2,"Sydsverige"
"Y_GE25","SE23",2013,5.5,"Västsverige"
"Y_GE25","SE3",2013,5.5,"Norra Sverige"
"Y_GE25","SE31",2013,6.2,"Norra Mellansverige"
"Y_GE25","SE32",2013,4.9,"Mellersta Norrland"
"Y_GE25","SE33",2013,4.9,"Övre Norrland"
"Y_GE25","SI",2013,9.2,"Slovenia"
"Y_GE25","SI0",2013,9.2,"Slovenija"
"Y_GE25","SI03",2013,10.2,"Vzhodna Slovenija"
"Y_GE25","SI04",2013,8.1,"Zahodna Slovenija"
"Y_GE25","SK",2013,12.5,"Slovakia"
"Y_GE25","SK0",2013,12.5,"Slovensko"
"Y_GE25","SK01",2013,5.6,"Bratislavský kraj"
"Y_GE25","SK02",2013,10.3,"Západné Slovensko"
"Y_GE25","SK03",2013,14.9,"Stredné Slovensko"
"Y_GE25","SK04",2013,16.4,"Východné Slovensko"
"Y_GE25","TR",2013,7.2,"Turkey"
"Y_GE25","TR1",2013,9.1,"Istanbul"
"Y_GE25","TR10",2013,9.1,"Istanbul"
"Y_GE25","TR2",2013,4.8,"Bati Marmara"
"Y_GE25","TR21",2013,5.3,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2013,4.2,"Balikesir, Çanakkale"
"Y_GE25","TR3",2013,7.7,"Ege"
"Y_GE25","TR31",2013,12.3,"Izmir"
"Y_GE25","TR32",2013,5,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2013,3.9,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2013,5.9,"Dogu Marmara"
"Y_GE25","TR41",2013,4.8,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2013,7.1,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2013,6,"Bati Anadolu"
"Y_GE25","TR51",2013,7.2,"Ankara"
"Y_GE25","TR52",2013,3,"Konya, Karaman"
"Y_GE25","TR6",2013,8.2,"Akdeniz"
"Y_GE25","TR61",2013,5.8,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2013,9.4,"Adana, Mersin"
"Y_GE25","TR63",2013,9.5,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2013,5.8,"Orta Anadolu"
"Y_GE25","TR71",2013,4.3,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2013,6.9,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2013,4.3,"Bati Karadeniz"
"Y_GE25","TR81",2013,4.8,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2013,4.3,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2013,4,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2013,4.4,"Dogu Karadeniz"
"Y_GE25","TR90",2013,4.4,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2013,4.9,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2013,5.1,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2013,4.7,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2013,5.6,"Ortadogu Anadolu"
"Y_GE25","TRB1",2013,4.3,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2013,7.1,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2013,11.2,"Güneydogu Anadolu"
"Y_GE25","TRC1",2013,5.3,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2013,14.6,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2013,16.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2013,5.4,"United Kingdom"
"Y_GE25","UKC",2013,7,"North East (UK)"
"Y_GE25","UKC1",2013,7.5,"Tees Valley and Durham"
"Y_GE25","UKC2",2013,6.7,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2013,6,"North West (UK)"
"Y_GE25","UKD1",2013,4,"Cumbria"
"Y_GE25","UKD3",2013,7.1,"Greater Manchester"
"Y_GE25","UKD4",2013,5,"Lancashire"
"Y_GE25","UKD6",2013,3.7,"Cheshire"
"Y_GE25","UKD7",2013,7.1,"Merseyside"
"Y_GE25","UKE",2013,6.1,"Yorkshire and The Humber"
"Y_GE25","UKE1",2013,6.2,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2013,3.1,"North Yorkshire"
"Y_GE25","UKE3",2013,7.2,"South Yorkshire"
"Y_GE25","UKE4",2013,6.4,"West Yorkshire"
"Y_GE25","UKF",2013,5.4,"East Midlands (UK)"
"Y_GE25","UKF1",2013,5,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2013,6.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2013,4.3,"Lincolnshire"
"Y_GE25","UKG",2013,6.5,"West Midlands (UK)"
"Y_GE25","UKG1",2013,3.7,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2013,4.7,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2013,9.2,"West Midlands"
"Y_GE25","UKH",2013,4.3,"East of England"
"Y_GE25","UKH1",2013,4.1,"East Anglia"
"Y_GE25","UKH2",2013,4.3,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2013,4.4,"Essex"
"Y_GE25","UKI",2013,6.5,"London"
"Y_GE25","UKI3",2013,6.1,"Inner London - West"
"Y_GE25","UKI4",2013,7.2,"Inner London - East"
"Y_GE25","UKI5",2013,7.2,"Outer London - East and North East"
"Y_GE25","UKI6",2013,4.5,"Outer London - South"
"Y_GE25","UKI7",2013,6.5,"Outer London - West and North West"
"Y_GE25","UKJ",2013,4,"South East (UK)"
"Y_GE25","UKJ1",2013,3.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2013,3.8,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2013,3.9,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2013,5.2,"Kent"
"Y_GE25","UKK",2013,4.3,"South West (UK)"
"Y_GE25","UKK1",2013,4.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2013,4,"Dorset and Somerset"
"Y_GE25","UKK3",2013,4.3,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2013,4.5,"Devon"
"Y_GE25","UKL",2013,5.2,"Wales"
"Y_GE25","UKL1",2013,5.5,"West Wales and The Valleys"
"Y_GE25","UKL2",2013,4.8,"East Wales"
"Y_GE25","UKM",2013,5.1,"Scotland"
"Y_GE25","UKM2",2013,4.5,"Eastern Scotland"
"Y_GE25","UKM3",2013,6.1,"South Western Scotland"
"Y_GE25","UKM5",2013,4,"North Eastern Scotland"
"Y_GE25","UKM6",2013,4.3,"Highlands and Islands"
"Y_GE25","UKN",2013,5.3,"Northern Ireland (UK)"
"Y_GE25","UKN0",2013,5.3,"Northern Ireland (UK)"
"Y15-24","AT",2012,9.4,"Austria"
"Y15-24","AT1",2012,13.4,"Ostösterreich"
"Y15-24","AT11",2012,NA,"Burgenland (AT)"
"Y15-24","AT12",2012,8.6,"Niederösterreich"
"Y15-24","AT13",2012,19.4,"Wien"
"Y15-24","AT2",2012,7.7,"Südösterreich"
"Y15-24","AT21",2012,12.1,"Kärnten"
"Y15-24","AT22",2012,5.8,"Steiermark"
"Y15-24","AT3",2012,6.6,"Westösterreich"
"Y15-24","AT31",2012,6.4,"Oberösterreich"
"Y15-24","AT32",2012,NA,"Salzburg"
"Y15-24","AT33",2012,6.4,"Tirol"
"Y15-24","AT34",2012,NA,"Vorarlberg"
"Y15-24","BE",2012,19.8,"Belgium"
"Y15-24","BE1",2012,36.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2012,36.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2012,12.8,"Vlaams Gewest"
"Y15-24","BE21",2012,11.7,"Prov. Antwerpen"
"Y15-24","BE22",2012,18.6,"Prov. Limburg (BE)"
"Y15-24","BE23",2012,11.8,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2012,15.1,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2012,9.9,"Prov. West-Vlaanderen"
"Y15-24","BE3",2012,27.1,"Région wallonne"
"Y15-24","BE31",2012,24.4,"Prov. Brabant Wallon"
"Y15-24","BE32",2012,32,"Prov. Hainaut"
"Y15-24","BE33",2012,25.8,"Prov. Liège"
"Y15-24","BE34",2012,23.1,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2012,21,"Prov. Namur"
"Y15-24","BG",2012,28.1,"Bulgaria"
"Y15-24","BG3",2012,33.6,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2012,30,"Severozapaden"
"Y15-24","BG32",2012,33.7,"Severen tsentralen"
"Y15-24","BG33",2012,36.1,"Severoiztochen"
"Y15-24","BG34",2012,33.4,"Yugoiztochen"
"Y15-24","BG4",2012,22.9,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2012,17.3,"Yugozapaden"
"Y15-24","BG42",2012,33.4,"Yuzhen tsentralen"
"Y15-24","CH",2012,8.4,"Switzerland"
"Y15-24","CH0",2012,8.4,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2012,14.1,"Région lémanique"
"Y15-24","CH02",2012,7.9,"Espace Mittelland"
"Y15-24","CH03",2012,8.8,"Nordwestschweiz"
"Y15-24","CH04",2012,6.6,"Zürich"
"Y15-24","CH05",2012,5.6,"Ostschweiz"
"Y15-24","CH06",2012,4.7,"Zentralschweiz"
"Y15-24","CH07",2012,18.1,"Ticino"
"Y15-24","CY",2012,27.7,"Cyprus"
"Y15-24","CY0",2012,27.7,"Kypros"
"Y15-24","CY00",2012,27.7,"Kypros"
"Y15-24","CZ",2012,19.5,"Czech Republic"
"Y15-24","CZ0",2012,19.5,"Ceská republika"
"Y15-24","CZ01",2012,11.9,"Praha"
"Y15-24","CZ02",2012,13.3,"Strední Cechy"
"Y15-24","CZ03",2012,13.2,"Jihozápad"
"Y15-24","CZ04",2012,28.2,"Severozápad"
"Y15-24","CZ05",2012,21.5,"Severovýchod"
"Y15-24","CZ06",2012,21.7,"Jihovýchod"
"Y15-24","CZ07",2012,21.2,"Strední Morava"
"Y15-24","CZ08",2012,20.9,"Moravskoslezsko"
"Y15-24","DE",2012,8,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2012,5.5,"Baden-Württemberg"
"Y15-24","DE11",2012,5.6,"Stuttgart"
"Y15-24","DE12",2012,6.8,"Karlsruhe"
"Y15-24","DE13",2012,4.8,"Freiburg"
"Y15-24","DE14",2012,4.4,"Tübingen"
"Y15-24","DE2",2012,5.3,"Bayern"
"Y15-24","DE21",2012,4.1,"Oberbayern"
"Y15-24","DE22",2012,5.9,"Niederbayern"
"Y15-24","DE23",2012,NA,"Oberpfalz"
"Y15-24","DE24",2012,NA,"Oberfranken"
"Y15-24","DE25",2012,6.8,"Mittelfranken"
"Y15-24","DE26",2012,NA,"Unterfranken"
"Y15-24","DE27",2012,5.3,"Schwaben"
"Y15-24","DE3",2012,14.9,"Berlin"
"Y15-24","DE30",2012,14.9,"Berlin"
"Y15-24","DE4",2012,13.3,"Brandenburg"
"Y15-24","DE40",2012,13.3,"Brandenburg"
"Y15-24","DE5",2012,NA,"Bremen"
"Y15-24","DE50",2012,NA,"Bremen"
"Y15-24","DE6",2012,7.2,"Hamburg"
"Y15-24","DE60",2012,7.2,"Hamburg"
"Y15-24","DE7",2012,7.8,"Hessen"
"Y15-24","DE71",2012,8.1,"Darmstadt"
"Y15-24","DE72",2012,NA,"Gießen"
"Y15-24","DE73",2012,NA,"Kassel"
"Y15-24","DE8",2012,12.9,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2012,12.9,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2012,7.9,"Niedersachsen"
"Y15-24","DE91",2012,9.7,"Braunschweig"
"Y15-24","DE92",2012,9.1,"Hannover"
"Y15-24","DE93",2012,6.5,"Lüneburg"
"Y15-24","DE94",2012,6.8,"Weser-Ems"
"Y15-24","DEA",2012,9.1,"Nordrhein-Westfalen"
"Y15-24","DEA1",2012,10,"Düsseldorf"
"Y15-24","DEA2",2012,8.2,"Köln"
"Y15-24","DEA3",2012,8.5,"Münster"
"Y15-24","DEA4",2012,8.8,"Detmold"
"Y15-24","DEA5",2012,9.4,"Arnsberg"
"Y15-24","DEB",2012,7,"Rheinland-Pfalz"
"Y15-24","DEB1",2012,5.7,"Koblenz"
"Y15-24","DEB2",2012,NA,"Trier"
"Y15-24","DEB3",2012,9.2,"Rheinhessen-Pfalz"
"Y15-24","DEC",2012,12.3,"Saarland"
"Y15-24","DEC0",2012,12.3,"Saarland"
"Y15-24","DED",2012,9.2,"Sachsen"
"Y15-24","DED2",2012,9.4,"Dresden"
"Y15-24","DED4",2012,9.1,"Chemnitz"
"Y15-24","DED5",2012,NA,"Leipzig"
"Y15-24","DEE",2012,13.4,"Sachsen-Anhalt"
"Y15-24","DEE0",2012,13.4,"Sachsen-Anhalt"
"Y15-24","DEF",2012,8.7,"Schleswig-Holstein"
"Y15-24","DEF0",2012,8.7,"Schleswig-Holstein"
"Y15-24","DEG",2012,9.1,"Thüringen"
"Y15-24","DEG0",2012,9.1,"Thüringen"
"Y15-24","DK",2012,14.1,"Denmark"
"Y15-24","DK0",2012,14.1,"Danmark"
"Y15-24","DK01",2012,14.1,"Hovedstaden"
"Y15-24","DK02",2012,15,"Sjælland"
"Y15-24","DK03",2012,14.6,"Syddanmark"
"Y15-24","DK04",2012,13.2,"Midtjylland"
"Y15-24","DK05",2012,14.4,"Nordjylland"
"Y15-24","EA17",2012,23.5,"Euro area (17 countries)"
"Y15-24","EA18",2012,23.6,"Euro area (18 countries)"
"Y15-24","EA19",2012,23.6,"Euro area (19 countries)"
"Y15-24","EE",2012,20.9,"Estonia"
"Y15-24","EE0",2012,20.9,"Eesti"
"Y15-24","EE00",2012,20.9,"Eesti"
"Y15-24","EL",2012,55.3,"Greece"
"Y15-24","EL3",2012,56,"Attiki"
"Y15-24","EL30",2012,56,"Attiki"
"Y15-24","EL4",2012,43.6,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2012,45.8,"Voreio Aigaio"
"Y15-24","EL42",2012,41,"Notio Aigaio"
"Y15-24","EL43",2012,44.1,"Kriti"
"Y15-24","EL5",2012,60,"Voreia Ellada"
"Y15-24","EL51",2012,53,"Anatoliki Makedonia, Thraki"
"Y15-24","EL52",2012,60.7,"Kentriki Makedonia"
"Y15-24","EL53",2012,72.3,"Dytiki Makedonia"
"Y15-24","EL54",2012,61.1,"Ipeiros"
"Y15-24","EL6",2012,55.1,"Kentriki Ellada"
"Y15-24","EL61",2012,53.7,"Thessalia"
"Y15-24","EL62",2012,23.9,"Ionia Nisia"
"Y15-24","EL63",2012,56.8,"Dytiki Ellada"
"Y15-24","EL64",2012,58.7,"Sterea Ellada"
"Y15-24","EL65",2012,62.3,"Peloponnisos"
"Y15-24","ES",2012,52.9,"Spain"
"Y15-24","ES1",2012,45.5,"Noroeste (ES)"
"Y15-24","ES11",2012,45.2,"Galicia"
"Y15-24","ES12",2012,48.9,"Principado de Asturias"
"Y15-24","ES13",2012,41.7,"Cantabria"
"Y15-24","ES2",2012,42.8,"Noreste (ES)"
"Y15-24","ES21",2012,42.7,"País Vasco"
"Y15-24","ES22",2012,40.1,"Comunidad Foral de Navarra"
"Y15-24","ES23",2012,50.1,"La Rioja"
"Y15-24","ES24",2012,42.4,"Aragón"
"Y15-24","ES3",2012,48.1,"Comunidad de Madrid"
"Y15-24","ES30",2012,48.1,"Comunidad de Madrid"
"Y15-24","ES4",2012,54,"Centro (ES)"
"Y15-24","ES41",2012,48.1,"Castilla y León"
"Y15-24","ES42",2012,54.5,"Castilla-la Mancha"
"Y15-24","ES43",2012,61.9,"Extremadura"
"Y15-24","ES5",2012,51.1,"Este (ES)"
"Y15-24","ES51",2012,50.4,"Cataluña"
"Y15-24","ES52",2012,52.9,"Comunidad Valenciana"
"Y15-24","ES53",2012,48.9,"Illes Balears"
"Y15-24","ES6",2012,60.3,"Sur (ES)"
"Y15-24","ES61",2012,61.9,"Andalucía"
"Y15-24","ES62",2012,50.4,"Región de Murcia"
"Y15-24","ES63",2012,70.4,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2012,60.1,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2012,62.3,"Canarias (ES)"
"Y15-24","ES70",2012,62.3,"Canarias (ES)"
"Y15-24","EU15",2012,22.7,"European Union (15 countries)"
"Y15-24","EU27",2012,23.2,"European Union (27 countries)"
"Y15-24","EU28",2012,23.3,"European Union (28 countries)"
"Y15-24","FI",2012,19,"Finland"
"Y15-24","FI1",2012,19,"Manner-Suomi"
"Y15-24","FI19",2012,21.3,"Länsi-Suomi"
"Y15-24","FI1B",2012,15.5,"Helsinki-Uusimaa"
"Y15-24","FI1C",2012,17.8,"Etelä-Suomi"
"Y15-24","FI1D",2012,22.2,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2012,NA,"Åland"
"Y15-24","FI20",2012,NA,"Åland"
"Y15-24","FR",2012,24.5,"France"
"Y15-24","FR1",2012,19.4,"Île de France"
"Y15-24","FR10",2012,19.4,"Île de France"
"Y15-24","FR2",2012,26.1,"Bassin Parisien"
"Y15-24","FR21",2012,25.4,"Champagne-Ardenne"
"Y15-24","FR22",2012,28.1,"Picardie"
"Y15-24","FR23",2012,26.7,"Haute-Normandie"
"Y15-24","FR24",2012,28.9,"Centre (FR)"
"Y15-24","FR25",2012,21.3,"Basse-Normandie"
"Y15-24","FR26",2012,23.6,"Bourgogne"
"Y15-24","FR3",2012,34.8,"Nord - Pas-de-Calais"
"Y15-24","FR30",2012,34.8,"Nord - Pas-de-Calais"
"Y15-24","FR4",2012,23.1,"Est (FR)"
"Y15-24","FR41",2012,24.4,"Lorraine"
"Y15-24","FR42",2012,22.9,"Alsace"
"Y15-24","FR43",2012,20.8,"Franche-Comté"
"Y15-24","FR5",2012,21.2,"Ouest (FR)"
"Y15-24","FR51",2012,22.2,"Pays de la Loire"
"Y15-24","FR52",2012,17.9,"Bretagne"
"Y15-24","FR53",2012,24.1,"Poitou-Charentes"
"Y15-24","FR6",2012,20.9,"Sud-Ouest (FR)"
"Y15-24","FR61",2012,24.7,"Aquitaine"
"Y15-24","FR62",2012,17.7,"Midi-Pyrénées"
"Y15-24","FR63",2012,NA,"Limousin"
"Y15-24","FR7",2012,20.9,"Centre-Est (FR)"
"Y15-24","FR71",2012,19.4,"Rhône-Alpes"
"Y15-24","FR72",2012,27.6,"Auvergne"
"Y15-24","FR8",2012,28.1,"Méditerranée"
"Y15-24","FR81",2012,38.2,"Languedoc-Roussillon"
"Y15-24","FR82",2012,22.2,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2012,NA,"Corse"
"Y15-24","FRA",2012,53.9,"Départements d'outre-mer"
"Y15-24","FRA1",2012,53,"Guadeloupe"
"Y15-24","FRA2",2012,56.7,"Martinique"
"Y15-24","FRA3",2012,49.5,"Guyane"
"Y15-24","FRA4",2012,54.2,"La Réunion"
"Y15-24","HR",2012,42.1,"Croatia"
"Y15-24","HR0",2012,42.1,"Hrvatska"
"Y15-24","HR03",2012,36.8,"Jadranska Hrvatska"
"Y15-24","HR04",2012,44.4,"Kontinentalna Hrvatska"
"Y15-24","HU",2012,28.2,"Hungary"
"Y15-24","HU1",2012,23.8,"Közép-Magyarország"
"Y15-24","HU10",2012,23.8,"Közép-Magyarország"
"Y15-24","HU2",2012,24.2,"Dunántúl"
"Y15-24","HU21",2012,24.2,"Közép-Dunántúl"
"Y15-24","HU22",2012,20.6,"Nyugat-Dunántúl"
"Y15-24","HU23",2012,29.1,"Dél-Dunántúl"
"Y15-24","HU3",2012,33.9,"Alföld és Észak"
"Y15-24","HU31",2012,38.4,"Észak-Magyarország"
"Y15-24","HU32",2012,35.6,"Észak-Alföld"
"Y15-24","HU33",2012,27.4,"Dél-Alföld"
"Y15-24","IE",2012,30.4,"Ireland"
"Y15-24","IE0",2012,30.4,"Éire/Ireland"
"Y15-24","IE01",2012,33.8,"Border, Midland and Western"
"Y15-24","IE02",2012,29.2,"Southern and Eastern"
"Y15-24","IS",2012,13.5,"Iceland"
"Y15-24","IS0",2012,13.5,"Ísland"
"Y15-24","IS00",2012,13.5,"Ísland"
"Y15-24","IT",2012,35.3,"Italy"
"Y15-24","ITC",2012,28.4,"Nord-Ovest"
"Y15-24","ITC1",2012,32.1,"Piemonte"
"Y15-24","ITC2",2012,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2012,30.2,"Liguria"
"Y15-24","ITC4",2012,26.5,"Lombardia"
"Y15-24","ITF",2012,45.5,"Sud"
"Y15-24","ITF1",2012,34,"Abruzzo"
"Y15-24","ITF2",2012,41.5,"Molise"
"Y15-24","ITF3",2012,48.4,"Campania"
"Y15-24","ITF4",2012,41.6,"Puglia"
"Y15-24","ITF5",2012,49.9,"Basilicata"
"Y15-24","ITF6",2012,53.9,"Calabria"
"Y15-24","ITG",2012,50.3,"Isole"
"Y15-24","ITG1",2012,51.2,"Sicilia"
"Y15-24","ITG2",2012,47.5,"Sardegna"
"Y15-24","ITH",2012,24,"Nord-Est"
"Y15-24","ITH1",2012,11.3,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2012,20.8,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2012,23.3,"Veneto"
"Y15-24","ITH4",2012,29.7,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2012,26.7,"Emilia-Romagna"
"Y15-24","ITI",2012,34.7,"Centro (IT)"
"Y15-24","ITI1",2012,29.4,"Toscana"
"Y15-24","ITI2",2012,34.6,"Umbria"
"Y15-24","ITI3",2012,28.6,"Marche"
"Y15-24","ITI4",2012,40,"Lazio"
"Y15-24","LT",2012,26.7,"Lithuania"
"Y15-24","LT0",2012,26.7,"Lietuva"
"Y15-24","LT00",2012,26.7,"Lietuva"
"Y15-24","LU",2012,18.8,"Luxembourg"
"Y15-24","LU0",2012,18.8,"Luxembourg"
"Y15-24","LU00",2012,18.8,"Luxembourg"
"Y15-24","LV",2012,28.5,"Latvia"
"Y15-24","LV0",2012,28.5,"Latvija"
"Y15-24","LV00",2012,28.5,"Latvija"
"Y15-24","MK",2012,53.9,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2012,53.9,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2012,53.9,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2012,14.1,"Malta"
"Y15-24","MT0",2012,14.1,"Malta"
"Y15-24","MT00",2012,14.1,"Malta"
"Y15-24","NL",2012,11.7,"Netherlands"
"Y15-24","NL1",2012,13,"Noord-Nederland"
"Y15-24","NL11",2012,14.4,"Groningen"
"Y15-24","NL12",2012,12.3,"Friesland (NL)"
"Y15-24","NL13",2012,12,"Drenthe"
"Y15-24","NL2",2012,11.4,"Oost-Nederland"
"Y15-24","NL21",2012,11.4,"Overijssel"
"Y15-24","NL22",2012,10.7,"Gelderland"
"Y15-24","NL23",2012,14.4,"Flevoland"
"Y15-24","NL3",2012,11.9,"West-Nederland"
"Y15-24","NL31",2012,10.4,"Utrecht"
"Y15-24","NL32",2012,10.8,"Noord-Holland"
"Y15-24","NL33",2012,13.7,"Zuid-Holland"
"Y15-24","NL34",2012,7.1,"Zeeland"
"Y15-24","NL4",2012,11,"Zuid-Nederland"
"Y15-24","NL41",2012,11.1,"Noord-Brabant"
"Y15-24","NL42",2012,10.9,"Limburg (NL)"
"Y15-24","NO",2012,8.5,"Norway"
"Y15-24","NO0",2012,8.5,"Norge"
"Y15-24","NO01",2012,9,"Oslo og Akershus"
"Y15-24","NO02",2012,6.5,"Hedmark og Oppland"
"Y15-24","NO03",2012,9.7,"Sør-Østlandet"
"Y15-24","NO04",2012,6.7,"Agder og Rogaland"
"Y15-24","NO05",2012,8.4,"Vestlandet"
"Y15-24","NO06",2012,8.8,"Trøndelag"
"Y15-24","NO07",2012,8.9,"Nord-Norge"
"Y15-24","PL",2012,26.5,"Poland"
"Y15-24","PL1",2012,22.3,"Region Centralny"
"Y15-24","PL11",2012,28.3,"Lódzkie"
"Y15-24","PL12",2012,19.4,"Mazowieckie"
"Y15-24","PL2",2012,24.7,"Region Poludniowy"
"Y15-24","PL21",2012,27.7,"Malopolskie"
"Y15-24","PL22",2012,22.3,"Slaskie"
"Y15-24","PL3",2012,32.9,"Region Wschodni"
"Y15-24","PL31",2012,30.9,"Lubelskie"
"Y15-24","PL32",2012,40.8,"Podkarpackie"
"Y15-24","PL33",2012,31.2,"Swietokrzyskie"
"Y15-24","PL34",2012,24.3,"Podlaskie"
"Y15-24","PL4",2012,25.2,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2012,22.9,"Wielkopolskie"
"Y15-24","PL42",2012,31.6,"Zachodniopomorskie"
"Y15-24","PL43",2012,26.4,"Lubuskie"
"Y15-24","PL5",2012,28,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2012,29.8,"Dolnoslaskie"
"Y15-24","PL52",2012,22.7,"Opolskie"
"Y15-24","PL6",2012,27.7,"Region Pólnocny"
"Y15-24","PL61",2012,30.5,"Kujawsko-Pomorskie"
"Y15-24","PL62",2012,29.3,"Warminsko-Mazurskie"
"Y15-24","PL63",2012,24.1,"Pomorskie"
"Y15-24","PT",2012,37.9,"Portugal"
"Y15-24","PT1",2012,37.5,"Continente"
"Y15-24","PT11",2012,33,"Norte"
"Y15-24","PT15",2012,40.5,"Algarve"
"Y15-24","PT16",2012,36.6,"Centro (PT)"
"Y15-24","PT17",2012,43.5,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2012,45,"Alentejo"
"Y15-24","PT2",2012,38.9,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2012,38.9,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2012,50.2,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2012,50.2,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2012,22.6,"Romania"
"Y15-24","RO1",2012,23.5,"Macroregiunea unu"
"Y15-24","RO11",2012,16.2,"Nord-Vest"
"Y15-24","RO12",2012,31.9,"Centru"
"Y15-24","RO2",2012,19.5,"Macroregiunea doi"
"Y15-24","RO21",2012,12.5,"Nord-Est"
"Y15-24","RO22",2012,30,"Sud-Est"
"Y15-24","RO3",2012,26.9,"Macroregiunea trei"
"Y15-24","RO31",2012,30,"Sud - Muntenia"
"Y15-24","RO32",2012,21.8,"Bucuresti - Ilfov"
"Y15-24","RO4",2012,19.9,"Macroregiunea patru"
"Y15-24","RO41",2012,19.6,"Sud-Vest Oltenia"
"Y15-24","RO42",2012,20.2,"Vest"
"Y15-24","SE",2012,23.6,"Sweden"
"Y15-24","SE1",2012,22.8,"Östra Sverige"
"Y15-24","SE11",2012,21.3,"Stockholm"
"Y15-24","SE12",2012,24.7,"Östra Mellansverige"
"Y15-24","SE2",2012,23.8,"Södra Sverige"
"Y15-24","SE21",2012,22.1,"Småland med öarna"
"Y15-24","SE22",2012,26.3,"Sydsverige"
"Y15-24","SE23",2012,22.8,"Västsverige"
"Y15-24","SE3",2012,25.1,"Norra Sverige"
"Y15-24","SE31",2012,25.2,"Norra Mellansverige"
"Y15-24","SE32",2012,26.4,"Mellersta Norrland"
"Y15-24","SE33",2012,24,"Övre Norrland"
"Y15-24","SI",2012,20.6,"Slovenia"
"Y15-24","SI0",2012,20.6,"Slovenija"
"Y15-24","SI03",2012,21.9,"Vzhodna Slovenija"
"Y15-24","SI04",2012,19,"Zahodna Slovenija"
"Y15-24","SK",2012,34,"Slovakia"
"Y15-24","SK0",2012,34,"Slovensko"
"Y15-24","SK01",2012,17.5,"Bratislavský kraj"
"Y15-24","SK02",2012,25.3,"Západné Slovensko"
"Y15-24","SK03",2012,38.8,"Stredné Slovensko"
"Y15-24","SK04",2012,43,"Východné Slovensko"
"Y15-24","TR",2012,15.7,"Turkey"
"Y15-24","TR1",2012,19.2,"Istanbul"
"Y15-24","TR10",2012,19.2,"Istanbul"
"Y15-24","TR2",2012,14.3,"Bati Marmara"
"Y15-24","TR21",2012,15.4,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2012,12.8,"Balikesir, Çanakkale"
"Y15-24","TR3",2012,16.2,"Ege"
"Y15-24","TR31",2012,23.6,"Izmir"
"Y15-24","TR32",2012,12.4,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2012,9.4,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2012,14.9,"Dogu Marmara"
"Y15-24","TR41",2012,12.1,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2012,17.7,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2012,16.5,"Bati Anadolu"
"Y15-24","TR51",2012,20.2,"Ankara"
"Y15-24","TR52",2012,10.4,"Konya, Karaman"
"Y15-24","TR6",2012,15.3,"Akdeniz"
"Y15-24","TR61",2012,13.5,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2012,15.2,"Adana, Mersin"
"Y15-24","TR63",2012,17.4,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2012,13.2,"Orta Anadolu"
"Y15-24","TR71",2012,15.8,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2012,11.8,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2012,10.6,"Bati Karadeniz"
"Y15-24","TR81",2012,16.2,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2012,9.1,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2012,8.6,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2012,19.3,"Dogu Karadeniz"
"Y15-24","TR90",2012,19.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2012,10.3,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2012,10.1,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2012,10.4,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2012,12.4,"Ortadogu Anadolu"
"Y15-24","TRB1",2012,13.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2012,11.5,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2012,16.2,"Güneydogu Anadolu"
"Y15-24","TRC1",2012,14.6,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2012,7.8,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2012,28.7,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2012,21.2,"United Kingdom"
"Y15-24","UKC",2012,24.7,"North East (UK)"
"Y15-24","UKC1",2012,33,"Tees Valley and Durham"
"Y15-24","UKC2",2012,19.2,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2012,23.4,"North West (UK)"
"Y15-24","UKD1",2012,15.5,"Cumbria"
"Y15-24","UKD3",2012,24.3,"Greater Manchester"
"Y15-24","UKD4",2012,24,"Lancashire"
"Y15-24","UKD6",2012,18.7,"Cheshire"
"Y15-24","UKD7",2012,25.5,"Merseyside"
"Y15-24","UKE",2012,22.9,"Yorkshire and The Humber"
"Y15-24","UKE1",2012,22,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2012,18.7,"North Yorkshire"
"Y15-24","UKE3",2012,21.4,"South Yorkshire"
"Y15-24","UKE4",2012,25.4,"West Yorkshire"
"Y15-24","UKF",2012,20.1,"East Midlands (UK)"
"Y15-24","UKF1",2012,22.3,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2012,17.2,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2012,20.3,"Lincolnshire"
"Y15-24","UKG",2012,23.3,"West Midlands (UK)"
"Y15-24","UKG1",2012,17.7,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2012,18.9,"Shropshire and Staffordshire"
"Y15-24","UKG3",2012,28,"West Midlands"
"Y15-24","UKH",2012,17.8,"East of England"
"Y15-24","UKH1",2012,17.3,"East Anglia"
"Y15-24","UKH2",2012,14.4,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2012,21.6,"Essex"
"Y15-24","UKI",2012,24.8,"London"
"Y15-24","UKI3",2012,21.7,"Inner London - West"
"Y15-24","UKI4",2012,27.7,"Inner London - East"
"Y15-24","UKI5",2012,25.5,"Outer London - East and North East"
"Y15-24","UKI6",2012,23.2,"Outer London - South"
"Y15-24","UKI7",2012,22.6,"Outer London - West and North West"
"Y15-24","UKJ",2012,17.9,"South East (UK)"
"Y15-24","UKJ1",2012,15.4,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2012,18,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2012,15.6,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2012,23.5,"Kent"
"Y15-24","UKK",2012,16,"South West (UK)"
"Y15-24","UKK1",2012,17,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2012,12.1,"Dorset and Somerset"
"Y15-24","UKK3",2012,14.6,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2012,18.7,"Devon"
"Y15-24","UKL",2012,24.2,"Wales"
"Y15-24","UKL1",2012,23.8,"West Wales and The Valleys"
"Y15-24","UKL2",2012,24.6,"East Wales"
"Y15-24","UKM",2012,21.6,"Scotland"
"Y15-24","UKM2",2012,20.5,"Eastern Scotland"
"Y15-24","UKM3",2012,24.7,"South Western Scotland"
"Y15-24","UKM5",2012,11.7,"North Eastern Scotland"
"Y15-24","UKM6",2012,24.6,"Highlands and Islands"
"Y15-24","UKN",2012,19.5,"Northern Ireland (UK)"
"Y15-24","UKN0",2012,19.5,"Northern Ireland (UK)"
"Y20-64","AT",2012,4.7,"Austria"
"Y20-64","AT1",2012,6.3,"Ostösterreich"
"Y20-64","AT11",2012,4.5,"Burgenland (AT)"
"Y20-64","AT12",2012,4.3,"Niederösterreich"
"Y20-64","AT13",2012,8.5,"Wien"
"Y20-64","AT2",2012,4.2,"Südösterreich"
"Y20-64","AT21",2012,4.8,"Kärnten"
"Y20-64","AT22",2012,3.9,"Steiermark"
"Y20-64","AT3",2012,3,"Westösterreich"
"Y20-64","AT31",2012,3.2,"Oberösterreich"
"Y20-64","AT32",2012,2.7,"Salzburg"
"Y20-64","AT33",2012,2.4,"Tirol"
"Y20-64","AT34",2012,3.7,"Vorarlberg"
"Y20-64","BE",2012,7.4,"Belgium"
"Y20-64","BE1",2012,17.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2012,17.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2012,4.3,"Vlaams Gewest"
"Y20-64","BE21",2012,5.1,"Prov. Antwerpen"
"Y20-64","BE22",2012,4.4,"Prov. Limburg (BE)"
"Y20-64","BE23",2012,4,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2012,4.3,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2012,3.7,"Prov. West-Vlaanderen"
"Y20-64","BE3",2012,9.8,"Région wallonne"
"Y20-64","BE31",2012,6.8,"Prov. Brabant Wallon"
"Y20-64","BE32",2012,11.9,"Prov. Hainaut"
"Y20-64","BE33",2012,10.5,"Prov. Liège"
"Y20-64","BE34",2012,7.4,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2012,7.2,"Prov. Namur"
"Y20-64","BG",2012,12,"Bulgaria"
"Y20-64","BG3",2012,13.9,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2012,11.7,"Severozapaden"
"Y20-64","BG32",2012,14,"Severen tsentralen"
"Y20-64","BG33",2012,17.9,"Severoiztochen"
"Y20-64","BG34",2012,11.6,"Yugoiztochen"
"Y20-64","BG4",2012,10.2,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2012,8.1,"Yugozapaden"
"Y20-64","BG42",2012,13.6,"Yuzhen tsentralen"
"Y20-64","CH",2012,4.1,"Switzerland"
"Y20-64","CH0",2012,4.1,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2012,6.4,"Région lémanique"
"Y20-64","CH02",2012,3.4,"Espace Mittelland"
"Y20-64","CH03",2012,4.1,"Nordwestschweiz"
"Y20-64","CH04",2012,3.5,"Zürich"
"Y20-64","CH05",2012,3.3,"Ostschweiz"
"Y20-64","CH06",2012,2.6,"Zentralschweiz"
"Y20-64","CH07",2012,7,"Ticino"
"Y20-64","CY",2012,11.8,"Cyprus"
"Y20-64","CY0",2012,11.8,"Kypros"
"Y20-64","CY00",2012,11.8,"Kypros"
"Y20-64","CZ",2012,6.8,"Czech Republic"
"Y20-64","CZ0",2012,6.8,"Ceská republika"
"Y20-64","CZ01",2012,3,"Praha"
"Y20-64","CZ02",2012,4.6,"Strední Cechy"
"Y20-64","CZ03",2012,5.1,"Jihozápad"
"Y20-64","CZ04",2012,10.2,"Severozápad"
"Y20-64","CZ05",2012,7.6,"Severovýchod"
"Y20-64","CZ06",2012,7.4,"Jihovýchod"
"Y20-64","CZ07",2012,7.4,"Strední Morava"
"Y20-64","CZ08",2012,9.3,"Moravskoslezsko"
"Y20-64","DE",2012,5.4,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2012,3.3,"Baden-Württemberg"
"Y20-64","DE11",2012,3.4,"Stuttgart"
"Y20-64","DE12",2012,4,"Karlsruhe"
"Y20-64","DE13",2012,2.8,"Freiburg"
"Y20-64","DE14",2012,2.6,"Tübingen"
"Y20-64","DE2",2012,3,"Bayern"
"Y20-64","DE21",2012,2.7,"Oberbayern"
"Y20-64","DE22",2012,3.2,"Niederbayern"
"Y20-64","DE23",2012,3.1,"Oberpfalz"
"Y20-64","DE24",2012,3.1,"Oberfranken"
"Y20-64","DE25",2012,3.4,"Mittelfranken"
"Y20-64","DE26",2012,3.3,"Unterfranken"
"Y20-64","DE27",2012,3.1,"Schwaben"
"Y20-64","DE3",2012,10.4,"Berlin"
"Y20-64","DE30",2012,10.4,"Berlin"
"Y20-64","DE4",2012,8.1,"Brandenburg"
"Y20-64","DE40",2012,8.1,"Brandenburg"
"Y20-64","DE5",2012,6.4,"Bremen"
"Y20-64","DE50",2012,6.4,"Bremen"
"Y20-64","DE6",2012,5.4,"Hamburg"
"Y20-64","DE60",2012,5.4,"Hamburg"
"Y20-64","DE7",2012,4.7,"Hessen"
"Y20-64","DE71",2012,4.7,"Darmstadt"
"Y20-64","DE72",2012,5,"Gießen"
"Y20-64","DE73",2012,4.5,"Kassel"
"Y20-64","DE8",2012,10.8,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2012,10.8,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2012,4.8,"Niedersachsen"
"Y20-64","DE91",2012,5.5,"Braunschweig"
"Y20-64","DE92",2012,5.4,"Hannover"
"Y20-64","DE93",2012,4.3,"Lüneburg"
"Y20-64","DE94",2012,4.2,"Weser-Ems"
"Y20-64","DEA",2012,5.8,"Nordrhein-Westfalen"
"Y20-64","DEA1",2012,6.4,"Düsseldorf"
"Y20-64","DEA2",2012,5.3,"Köln"
"Y20-64","DEA3",2012,4.9,"Münster"
"Y20-64","DEA4",2012,4.7,"Detmold"
"Y20-64","DEA5",2012,6.6,"Arnsberg"
"Y20-64","DEB",2012,3.9,"Rheinland-Pfalz"
"Y20-64","DEB1",2012,3.9,"Koblenz"
"Y20-64","DEB2",2012,2.7,"Trier"
"Y20-64","DEB3",2012,4.2,"Rheinhessen-Pfalz"
"Y20-64","DEC",2012,6.1,"Saarland"
"Y20-64","DEC0",2012,6.1,"Saarland"
"Y20-64","DED",2012,8.3,"Sachsen"
"Y20-64","DED2",2012,7.7,"Dresden"
"Y20-64","DED4",2012,8.1,"Chemnitz"
"Y20-64","DED5",2012,9.7,"Leipzig"
"Y20-64","DEE",2012,9.6,"Sachsen-Anhalt"
"Y20-64","DEE0",2012,9.6,"Sachsen-Anhalt"
"Y20-64","DEF",2012,4.9,"Schleswig-Holstein"
"Y20-64","DEF0",2012,4.9,"Schleswig-Holstein"
"Y20-64","DEG",2012,7.3,"Thüringen"
"Y20-64","DEG0",2012,7.3,"Thüringen"
"Y20-64","DK",2012,7,"Denmark"
"Y20-64","DK0",2012,7,"Danmark"
"Y20-64","DK01",2012,7.7,"Hovedstaden"
"Y20-64","DK02",2012,5.8,"Sjælland"
"Y20-64","DK03",2012,7.3,"Syddanmark"
"Y20-64","DK04",2012,6.4,"Midtjylland"
"Y20-64","DK05",2012,7.5,"Nordjylland"
"Y20-64","EA17",2012,11.1,"Euro area (17 countries)"
"Y20-64","EA18",2012,11.2,"Euro area (18 countries)"
"Y20-64","EA19",2012,11.2,"Euro area (19 countries)"
"Y20-64","EE",2012,10,"Estonia"
"Y20-64","EE0",2012,10,"Eesti"
"Y20-64","EE00",2012,10,"Eesti"
"Y20-64","EL",2012,24.3,"Greece"
"Y20-64","EL3",2012,25.6,"Attiki"
"Y20-64","EL30",2012,25.6,"Attiki"
"Y20-64","EL4",2012,20,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2012,20.9,"Voreio Aigaio"
"Y20-64","EL42",2012,15.1,"Notio Aigaio"
"Y20-64","EL43",2012,22.3,"Kriti"
"Y20-64","EL5",2012,25.3,"Voreia Ellada"
"Y20-64","EL51",2012,22.6,"Anatoliki Makedonia, Thraki"
"Y20-64","EL52",2012,26.1,"Kentriki Makedonia"
"Y20-64","EL53",2012,29.6,"Dytiki Makedonia"
"Y20-64","EL54",2012,22.5,"Ipeiros"
"Y20-64","EL6",2012,23,"Kentriki Ellada"
"Y20-64","EL61",2012,22.8,"Thessalia"
"Y20-64","EL62",2012,14.9,"Ionia Nisia"
"Y20-64","EL63",2012,25.4,"Dytiki Ellada"
"Y20-64","EL64",2012,27.5,"Sterea Ellada"
"Y20-64","EL65",2012,19.1,"Peloponnisos"
"Y20-64","ES",2012,24.3,"Spain"
"Y20-64","ES1",2012,20.4,"Noroeste (ES)"
"Y20-64","ES11",2012,20.4,"Galicia"
"Y20-64","ES12",2012,21.8,"Principado de Asturias"
"Y20-64","ES13",2012,17.7,"Cantabria"
"Y20-64","ES2",2012,16.6,"Noreste (ES)"
"Y20-64","ES21",2012,15.4,"País Vasco"
"Y20-64","ES22",2012,15.9,"Comunidad Foral de Navarra"
"Y20-64","ES23",2012,20.1,"La Rioja"
"Y20-64","ES24",2012,18.2,"Aragón"
"Y20-64","ES3",2012,18.1,"Comunidad de Madrid"
"Y20-64","ES30",2012,18.1,"Comunidad de Madrid"
"Y20-64","ES4",2012,25,"Centro (ES)"
"Y20-64","ES41",2012,19.4,"Castilla y León"
"Y20-64","ES42",2012,27.9,"Castilla-la Mancha"
"Y20-64","ES43",2012,32.4,"Extremadura"
"Y20-64","ES5",2012,23.7,"Este (ES)"
"Y20-64","ES51",2012,21.9,"Cataluña"
"Y20-64","ES52",2012,26.7,"Comunidad Valenciana"
"Y20-64","ES53",2012,22.6,"Illes Balears"
"Y20-64","ES6",2012,32.7,"Sur (ES)"
"Y20-64","ES61",2012,33.7,"Andalucía"
"Y20-64","ES62",2012,27,"Región de Murcia"
"Y20-64","ES63",2012,36.1,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2012,26,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2012,32.2,"Canarias (ES)"
"Y20-64","ES70",2012,32.2,"Canarias (ES)"
"Y20-64","EU15",2012,10.3,"European Union (15 countries)"
"Y20-64","EU27",2012,10.1,"European Union (27 countries)"
"Y20-64","EU28",2012,10.2,"European Union (28 countries)"
"Y20-64","FI",2012,7,"Finland"
"Y20-64","FI1",2012,7,"Manner-Suomi"
"Y20-64","FI19",2012,7.4,"Länsi-Suomi"
"Y20-64","FI1B",2012,5.6,"Helsinki-Uusimaa"
"Y20-64","FI1C",2012,6.7,"Etelä-Suomi"
"Y20-64","FI1D",2012,8.8,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2012,NA,"Åland"
"Y20-64","FI20",2012,NA,"Åland"
"Y20-64","FR",2012,9.4,"France"
"Y20-64","FR1",2012,7.9,"Île de France"
"Y20-64","FR10",2012,7.9,"Île de France"
"Y20-64","FR2",2012,9.7,"Bassin Parisien"
"Y20-64","FR21",2012,10.2,"Champagne-Ardenne"
"Y20-64","FR22",2012,10.1,"Picardie"
"Y20-64","FR23",2012,10.4,"Haute-Normandie"
"Y20-64","FR24",2012,10.3,"Centre (FR)"
"Y20-64","FR25",2012,8.4,"Basse-Normandie"
"Y20-64","FR26",2012,8.5,"Bourgogne"
"Y20-64","FR3",2012,12.4,"Nord - Pas-de-Calais"
"Y20-64","FR30",2012,12.4,"Nord - Pas-de-Calais"
"Y20-64","FR4",2012,9.5,"Est (FR)"
"Y20-64","FR41",2012,11.3,"Lorraine"
"Y20-64","FR42",2012,7.9,"Alsace"
"Y20-64","FR43",2012,8.7,"Franche-Comté"
"Y20-64","FR5",2012,7.8,"Ouest (FR)"
"Y20-64","FR51",2012,7.9,"Pays de la Loire"
"Y20-64","FR52",2012,7.7,"Bretagne"
"Y20-64","FR53",2012,7.9,"Poitou-Charentes"
"Y20-64","FR6",2012,8.5,"Sud-Ouest (FR)"
"Y20-64","FR61",2012,9.1,"Aquitaine"
"Y20-64","FR62",2012,8.2,"Midi-Pyrénées"
"Y20-64","FR63",2012,6.7,"Limousin"
"Y20-64","FR7",2012,8,"Centre-Est (FR)"
"Y20-64","FR71",2012,7.7,"Rhône-Alpes"
"Y20-64","FR72",2012,9.4,"Auvergne"
"Y20-64","FR8",2012,10.8,"Méditerranée"
"Y20-64","FR81",2012,14.2,"Languedoc-Roussillon"
"Y20-64","FR82",2012,9.3,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2012,7.3,"Corse"
"Y20-64","FRA",2012,24.4,"Départements d'outre-mer"
"Y20-64","FRA1",2012,22.7,"Guadeloupe"
"Y20-64","FRA2",2012,20.7,"Martinique"
"Y20-64","FRA3",2012,21.8,"Guyane"
"Y20-64","FRA4",2012,27.5,"La Réunion"
"Y20-64","HR",2012,15.5,"Croatia"
"Y20-64","HR0",2012,15.5,"Hrvatska"
"Y20-64","HR03",2012,14.2,"Jadranska Hrvatska"
"Y20-64","HR04",2012,16,"Kontinentalna Hrvatska"
"Y20-64","HU",2012,10.9,"Hungary"
"Y20-64","HU1",2012,9.4,"Közép-Magyarország"
"Y20-64","HU10",2012,9.4,"Közép-Magyarország"
"Y20-64","HU2",2012,9.6,"Dunántúl"
"Y20-64","HU21",2012,9.7,"Közép-Dunántúl"
"Y20-64","HU22",2012,7.4,"Nyugat-Dunántúl"
"Y20-64","HU23",2012,12,"Dél-Dunántúl"
"Y20-64","HU3",2012,13.1,"Alföld és Észak"
"Y20-64","HU31",2012,15.9,"Észak-Magyarország"
"Y20-64","HU32",2012,13.7,"Észak-Alföld"
"Y20-64","HU33",2012,10.2,"Dél-Alföld"
"Y20-64","IE",2012,14.4,"Ireland"
"Y20-64","IE0",2012,14.4,"Éire/Ireland"
"Y20-64","IE01",2012,16.2,"Border, Midland and Western"
"Y20-64","IE02",2012,13.8,"Southern and Eastern"
"Y20-64","IS",2012,5.3,"Iceland"
"Y20-64","IS0",2012,5.3,"Ísland"
"Y20-64","IS00",2012,5.3,"Ísland"
"Y20-64","IT",2012,10.3,"Italy"
"Y20-64","ITC",2012,7.6,"Nord-Ovest"
"Y20-64","ITC1",2012,8.9,"Piemonte"
"Y20-64","ITC2",2012,6.9,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2012,7.9,"Liguria"
"Y20-64","ITC4",2012,7.1,"Lombardia"
"Y20-64","ITF",2012,16.5,"Sud"
"Y20-64","ITF1",2012,10.5,"Abruzzo"
"Y20-64","ITF2",2012,11.8,"Molise"
"Y20-64","ITF3",2012,18.7,"Campania"
"Y20-64","ITF4",2012,15.2,"Puglia"
"Y20-64","ITF5",2012,14.3,"Basilicata"
"Y20-64","ITF6",2012,19,"Calabria"
"Y20-64","ITG",2012,17.2,"Isole"
"Y20-64","ITG1",2012,18,"Sicilia"
"Y20-64","ITG2",2012,15.2,"Sardegna"
"Y20-64","ITH",2012,6.3,"Nord-Est"
"Y20-64","ITH1",2012,3.8,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2012,5.8,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2012,6.2,"Veneto"
"Y20-64","ITH4",2012,6.6,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2012,6.8,"Emilia-Romagna"
"Y20-64","ITI",2012,9.2,"Centro (IT)"
"Y20-64","ITI1",2012,7.7,"Toscana"
"Y20-64","ITI2",2012,9,"Umbria"
"Y20-64","ITI3",2012,8.7,"Marche"
"Y20-64","ITI4",2012,10.4,"Lazio"
"Y20-64","LT",2012,13.5,"Lithuania"
"Y20-64","LT0",2012,13.5,"Lietuva"
"Y20-64","LT00",2012,13.5,"Lietuva"
"Y20-64","LU",2012,5,"Luxembourg"
"Y20-64","LU0",2012,5,"Luxembourg"
"Y20-64","LU00",2012,5,"Luxembourg"
"Y20-64","LV",2012,14.9,"Latvia"
"Y20-64","LV0",2012,14.9,"Latvija"
"Y20-64","LV00",2012,14.9,"Latvija"
"Y20-64","MK",2012,30.7,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2012,30.7,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2012,30.7,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2012,5.5,"Malta"
"Y20-64","MT0",2012,5.5,"Malta"
"Y20-64","MT00",2012,5.5,"Malta"
"Y20-64","NL",2012,5.2,"Netherlands"
"Y20-64","NL1",2012,6,"Noord-Nederland"
"Y20-64","NL11",2012,6.3,"Groningen"
"Y20-64","NL12",2012,5.7,"Friesland (NL)"
"Y20-64","NL13",2012,5.8,"Drenthe"
"Y20-64","NL2",2012,5,"Oost-Nederland"
"Y20-64","NL21",2012,5,"Overijssel"
"Y20-64","NL22",2012,4.7,"Gelderland"
"Y20-64","NL23",2012,6.5,"Flevoland"
"Y20-64","NL3",2012,5.3,"West-Nederland"
"Y20-64","NL31",2012,4.5,"Utrecht"
"Y20-64","NL32",2012,4.9,"Noord-Holland"
"Y20-64","NL33",2012,6.3,"Zuid-Holland"
"Y20-64","NL34",2012,3,"Zeeland"
"Y20-64","NL4",2012,4.7,"Zuid-Nederland"
"Y20-64","NL41",2012,4.7,"Noord-Brabant"
"Y20-64","NL42",2012,4.6,"Limburg (NL)"
"Y20-64","NO",2012,2.8,"Norway"
"Y20-64","NO0",2012,2.8,"Norge"
"Y20-64","NO01",2012,2.8,"Oslo og Akershus"
"Y20-64","NO02",2012,2.8,"Hedmark og Oppland"
"Y20-64","NO03",2012,3.2,"Sør-Østlandet"
"Y20-64","NO04",2012,2.4,"Agder og Rogaland"
"Y20-64","NO05",2012,2.5,"Vestlandet"
"Y20-64","NO06",2012,2.8,"Trøndelag"
"Y20-64","NO07",2012,3,"Nord-Norge"
"Y20-64","PL",2012,10,"Poland"
"Y20-64","PL1",2012,8.9,"Region Centralny"
"Y20-64","PL11",2012,10.9,"Lódzkie"
"Y20-64","PL12",2012,7.9,"Mazowieckie"
"Y20-64","PL2",2012,9.7,"Region Poludniowy"
"Y20-64","PL21",2012,10.3,"Malopolskie"
"Y20-64","PL22",2012,9.3,"Slaskie"
"Y20-64","PL3",2012,11.7,"Region Wschodni"
"Y20-64","PL31",2012,10.4,"Lubelskie"
"Y20-64","PL32",2012,13.3,"Podkarpackie"
"Y20-64","PL33",2012,13.3,"Swietokrzyskie"
"Y20-64","PL34",2012,9.2,"Podlaskie"
"Y20-64","PL4",2012,9,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2012,8.4,"Wielkopolskie"
"Y20-64","PL42",2012,10.7,"Zachodniopomorskie"
"Y20-64","PL43",2012,8.8,"Lubuskie"
"Y20-64","PL5",2012,10.5,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2012,10.9,"Dolnoslaskie"
"Y20-64","PL52",2012,9.3,"Opolskie"
"Y20-64","PL6",2012,10.6,"Region Pólnocny"
"Y20-64","PL61",2012,11.7,"Kujawsko-Pomorskie"
"Y20-64","PL62",2012,10.8,"Warminsko-Mazurskie"
"Y20-64","PL63",2012,9.4,"Pomorskie"
"Y20-64","PT",2012,15.8,"Portugal"
"Y20-64","PT1",2012,15.8,"Continente"
"Y20-64","PT11",2012,16.2,"Norte"
"Y20-64","PT15",2012,17.9,"Algarve"
"Y20-64","PT16",2012,12.2,"Centro (PT)"
"Y20-64","PT17",2012,17.5,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2012,16.2,"Alentejo"
"Y20-64","PT2",2012,14.9,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2012,14.9,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2012,17.3,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2012,17.3,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2012,6.7,"Romania"
"Y20-64","RO1",2012,6.6,"Macroregiunea unu"
"Y20-64","RO11",2012,4.5,"Nord-Vest"
"Y20-64","RO12",2012,9.1,"Centru"
"Y20-64","RO2",2012,6.4,"Macroregiunea doi"
"Y20-64","RO21",2012,4.3,"Nord-Est"
"Y20-64","RO22",2012,9.2,"Sud-Est"
"Y20-64","RO3",2012,8.1,"Macroregiunea trei"
"Y20-64","RO31",2012,9.5,"Sud - Muntenia"
"Y20-64","RO32",2012,6.4,"Bucuresti - Ilfov"
"Y20-64","RO4",2012,5.6,"Macroregiunea patru"
"Y20-64","RO41",2012,6.3,"Sud-Vest Oltenia"
"Y20-64","RO42",2012,4.8,"Vest"
"Y20-64","SE",2012,7.1,"Sweden"
"Y20-64","SE1",2012,6.5,"Östra Sverige"
"Y20-64","SE11",2012,5.8,"Stockholm"
"Y20-64","SE12",2012,7.6,"Östra Mellansverige"
"Y20-64","SE2",2012,7.4,"Södra Sverige"
"Y20-64","SE21",2012,6.6,"Småland med öarna"
"Y20-64","SE22",2012,8.5,"Sydsverige"
"Y20-64","SE23",2012,6.9,"Västsverige"
"Y20-64","SE3",2012,7.5,"Norra Sverige"
"Y20-64","SE31",2012,7.9,"Norra Mellansverige"
"Y20-64","SE32",2012,7.4,"Mellersta Norrland"
"Y20-64","SE33",2012,6.8,"Övre Norrland"
"Y20-64","SI",2012,8.9,"Slovenia"
"Y20-64","SI0",2012,8.9,"Slovenija"
"Y20-64","SI03",2012,10,"Vzhodna Slovenija"
"Y20-64","SI04",2012,7.6,"Zahodna Slovenija"
"Y20-64","SK",2012,13.6,"Slovakia"
"Y20-64","SK0",2012,13.6,"Slovensko"
"Y20-64","SK01",2012,5.6,"Bratislavský kraj"
"Y20-64","SK02",2012,11.1,"Západné Slovensko"
"Y20-64","SK03",2012,15.6,"Stredné Slovensko"
"Y20-64","SK04",2012,18.4,"Východné Slovensko"
"Y20-64","TR",2012,8,"Turkey"
"Y20-64","TR1",2012,10.4,"Istanbul"
"Y20-64","TR10",2012,10.4,"Istanbul"
"Y20-64","TR2",2012,5.3,"Bati Marmara"
"Y20-64","TR21",2012,6.1,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2012,4.4,"Balikesir, Çanakkale"
"Y20-64","TR3",2012,8.6,"Ege"
"Y20-64","TR31",2012,13,"Izmir"
"Y20-64","TR32",2012,6.8,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2012,4.1,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2012,7.4,"Dogu Marmara"
"Y20-64","TR41",2012,6.2,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2012,8.6,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2012,7.1,"Bati Anadolu"
"Y20-64","TR51",2012,8.1,"Ankara"
"Y20-64","TR52",2012,4.7,"Konya, Karaman"
"Y20-64","TR6",2012,8.3,"Akdeniz"
"Y20-64","TR61",2012,7.2,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2012,9,"Adana, Mersin"
"Y20-64","TR63",2012,8.7,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2012,6.9,"Orta Anadolu"
"Y20-64","TR71",2012,6,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2012,7.4,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2012,5.4,"Bati Karadeniz"
"Y20-64","TR81",2012,6.6,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2012,5,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2012,5,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2012,5.3,"Dogu Karadeniz"
"Y20-64","TR90",2012,5.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2012,5.8,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2012,5.5,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2012,6,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2012,6.6,"Ortadogu Anadolu"
"Y20-64","TRB1",2012,6,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2012,7.3,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2012,10.8,"Güneydogu Anadolu"
"Y20-64","TRC1",2012,10.7,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2012,6,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2012,17.6,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2012,6.9,"United Kingdom"
"Y20-64","UKC",2012,8.8,"North East (UK)"
"Y20-64","UKC1",2012,9.7,"Tees Valley and Durham"
"Y20-64","UKC2",2012,8.2,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2012,7.6,"North West (UK)"
"Y20-64","UKD1",2012,5.8,"Cumbria"
"Y20-64","UKD3",2012,8.6,"Greater Manchester"
"Y20-64","UKD4",2012,6.8,"Lancashire"
"Y20-64","UKD6",2012,5.6,"Cheshire"
"Y20-64","UKD7",2012,8.5,"Merseyside"
"Y20-64","UKE",2012,7.9,"Yorkshire and The Humber"
"Y20-64","UKE1",2012,8.7,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2012,4.3,"North Yorkshire"
"Y20-64","UKE3",2012,9.3,"South Yorkshire"
"Y20-64","UKE4",2012,8,"West Yorkshire"
"Y20-64","UKF",2012,6.7,"East Midlands (UK)"
"Y20-64","UKF1",2012,7.2,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2012,6,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2012,7.3,"Lincolnshire"
"Y20-64","UKG",2012,7.6,"West Midlands (UK)"
"Y20-64","UKG1",2012,4.4,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2012,5.6,"Shropshire and Staffordshire"
"Y20-64","UKG3",2012,10.4,"West Midlands"
"Y20-64","UKH",2012,5.7,"East of England"
"Y20-64","UKH1",2012,5.3,"East Anglia"
"Y20-64","UKH2",2012,5.7,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2012,6.4,"Essex"
"Y20-64","UKI",2012,8.2,"London"
"Y20-64","UKI3",2012,6.2,"Inner London - West"
"Y20-64","UKI4",2012,9.9,"Inner London - East"
"Y20-64","UKI5",2012,8.3,"Outer London - East and North East"
"Y20-64","UKI6",2012,6.3,"Outer London - South"
"Y20-64","UKI7",2012,8.6,"Outer London - West and North West"
"Y20-64","UKJ",2012,5.4,"South East (UK)"
"Y20-64","UKJ1",2012,4.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2012,4.8,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2012,5.5,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2012,7.1,"Kent"
"Y20-64","UKK",2012,5.1,"South West (UK)"
"Y20-64","UKK1",2012,5.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2012,4.3,"Dorset and Somerset"
"Y20-64","UKK3",2012,4.9,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2012,5.2,"Devon"
"Y20-64","UKL",2012,7.3,"Wales"
"Y20-64","UKL1",2012,8.3,"West Wales and The Valleys"
"Y20-64","UKL2",2012,5.8,"East Wales"
"Y20-64","UKM",2012,7,"Scotland"
"Y20-64","UKM2",2012,6.6,"Eastern Scotland"
"Y20-64","UKM3",2012,8.1,"South Western Scotland"
"Y20-64","UKM5",2012,4.3,"North Eastern Scotland"
"Y20-64","UKM6",2012,7.5,"Highlands and Islands"
"Y20-64","UKN",2012,7.2,"Northern Ireland (UK)"
"Y20-64","UKN0",2012,7.2,"Northern Ireland (UK)"
"Y_GE15","AT",2012,4.9,"Austria"
"Y_GE15","AT1",2012,6.6,"Ostösterreich"
"Y_GE15","AT11",2012,4.6,"Burgenland (AT)"
"Y_GE15","AT12",2012,4.6,"Niederösterreich"
"Y_GE15","AT13",2012,8.9,"Wien"
"Y_GE15","AT2",2012,4.3,"Südösterreich"
"Y_GE15","AT21",2012,5,"Kärnten"
"Y_GE15","AT22",2012,4,"Steiermark"
"Y_GE15","AT3",2012,3.2,"Westösterreich"
"Y_GE15","AT31",2012,3.3,"Oberösterreich"
"Y_GE15","AT32",2012,2.9,"Salzburg"
"Y_GE15","AT33",2012,2.8,"Tirol"
"Y_GE15","AT34",2012,4,"Vorarlberg"
"Y_GE15","BE",2012,7.5,"Belgium"
"Y_GE15","BE1",2012,17.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2012,17.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2012,4.5,"Vlaams Gewest"
"Y_GE15","BE21",2012,5.3,"Prov. Antwerpen"
"Y_GE15","BE22",2012,4.7,"Prov. Limburg (BE)"
"Y_GE15","BE23",2012,4.1,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2012,4.4,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2012,3.9,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2012,10,"Région wallonne"
"Y_GE15","BE31",2012,7,"Prov. Brabant Wallon"
"Y_GE15","BE32",2012,12.1,"Prov. Hainaut"
"Y_GE15","BE33",2012,10.7,"Prov. Liège"
"Y_GE15","BE34",2012,7.6,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2012,7.3,"Prov. Namur"
"Y_GE15","BG",2012,12.3,"Bulgaria"
"Y_GE15","BG3",2012,14.3,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2012,12.3,"Severozapaden"
"Y_GE15","BG32",2012,14.3,"Severen tsentralen"
"Y_GE15","BG33",2012,18.2,"Severoiztochen"
"Y_GE15","BG34",2012,11.9,"Yugoiztochen"
"Y_GE15","BG4",2012,10.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2012,8.2,"Yugozapaden"
"Y_GE15","BG42",2012,13.8,"Yuzhen tsentralen"
"Y_GE15","CH",2012,4.2,"Switzerland"
"Y_GE15","CH0",2012,4.2,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2012,6.6,"Région lémanique"
"Y_GE15","CH02",2012,3.5,"Espace Mittelland"
"Y_GE15","CH03",2012,4.1,"Nordwestschweiz"
"Y_GE15","CH04",2012,3.6,"Zürich"
"Y_GE15","CH05",2012,3.3,"Ostschweiz"
"Y_GE15","CH06",2012,2.7,"Zentralschweiz"
"Y_GE15","CH07",2012,6.9,"Ticino"
"Y_GE15","CY",2012,11.8,"Cyprus"
"Y_GE15","CY0",2012,11.8,"Kypros"
"Y_GE15","CY00",2012,11.8,"Kypros"
"Y_GE15","CZ",2012,7,"Czech Republic"
"Y_GE15","CZ0",2012,7,"Ceská republika"
"Y_GE15","CZ01",2012,3.1,"Praha"
"Y_GE15","CZ02",2012,4.6,"Strední Cechy"
"Y_GE15","CZ03",2012,5.3,"Jihozápad"
"Y_GE15","CZ04",2012,10.7,"Severozápad"
"Y_GE15","CZ05",2012,8,"Severovýchod"
"Y_GE15","CZ06",2012,7.6,"Jihovýchod"
"Y_GE15","CZ07",2012,7.5,"Strední Morava"
"Y_GE15","CZ08",2012,9.5,"Moravskoslezsko"
"Y_GE15","DE",2012,5.4,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2012,3.3,"Baden-Württemberg"
"Y_GE15","DE11",2012,3.4,"Stuttgart"
"Y_GE15","DE12",2012,4,"Karlsruhe"
"Y_GE15","DE13",2012,2.8,"Freiburg"
"Y_GE15","DE14",2012,2.7,"Tübingen"
"Y_GE15","DE2",2012,3.1,"Bayern"
"Y_GE15","DE21",2012,2.7,"Oberbayern"
"Y_GE15","DE22",2012,3.3,"Niederbayern"
"Y_GE15","DE23",2012,3.2,"Oberpfalz"
"Y_GE15","DE24",2012,3.3,"Oberfranken"
"Y_GE15","DE25",2012,3.7,"Mittelfranken"
"Y_GE15","DE26",2012,3.4,"Unterfranken"
"Y_GE15","DE27",2012,3.2,"Schwaben"
"Y_GE15","DE3",2012,10.4,"Berlin"
"Y_GE15","DE30",2012,10.4,"Berlin"
"Y_GE15","DE4",2012,8.2,"Brandenburg"
"Y_GE15","DE40",2012,8.2,"Brandenburg"
"Y_GE15","DE5",2012,6.6,"Bremen"
"Y_GE15","DE50",2012,6.6,"Bremen"
"Y_GE15","DE6",2012,5.3,"Hamburg"
"Y_GE15","DE60",2012,5.3,"Hamburg"
"Y_GE15","DE7",2012,4.7,"Hessen"
"Y_GE15","DE71",2012,4.8,"Darmstadt"
"Y_GE15","DE72",2012,5,"Gießen"
"Y_GE15","DE73",2012,4.5,"Kassel"
"Y_GE15","DE8",2012,10.8,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2012,10.8,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2012,4.9,"Niedersachsen"
"Y_GE15","DE91",2012,5.5,"Braunschweig"
"Y_GE15","DE92",2012,5.4,"Hannover"
"Y_GE15","DE93",2012,4.4,"Lüneburg"
"Y_GE15","DE94",2012,4.3,"Weser-Ems"
"Y_GE15","DEA",2012,5.8,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2012,6.5,"Düsseldorf"
"Y_GE15","DEA2",2012,5.4,"Köln"
"Y_GE15","DEA3",2012,4.9,"Münster"
"Y_GE15","DEA4",2012,4.7,"Detmold"
"Y_GE15","DEA5",2012,6.6,"Arnsberg"
"Y_GE15","DEB",2012,4,"Rheinland-Pfalz"
"Y_GE15","DEB1",2012,4,"Koblenz"
"Y_GE15","DEB2",2012,2.7,"Trier"
"Y_GE15","DEB3",2012,4.3,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2012,6.2,"Saarland"
"Y_GE15","DEC0",2012,6.2,"Saarland"
"Y_GE15","DED",2012,8.2,"Sachsen"
"Y_GE15","DED2",2012,7.5,"Dresden"
"Y_GE15","DED4",2012,7.9,"Chemnitz"
"Y_GE15","DED5",2012,9.5,"Leipzig"
"Y_GE15","DEE",2012,9.5,"Sachsen-Anhalt"
"Y_GE15","DEE0",2012,9.5,"Sachsen-Anhalt"
"Y_GE15","DEF",2012,5,"Schleswig-Holstein"
"Y_GE15","DEF0",2012,5,"Schleswig-Holstein"
"Y_GE15","DEG",2012,7.2,"Thüringen"
"Y_GE15","DEG0",2012,7.2,"Thüringen"
"Y_GE15","DK",2012,7.5,"Denmark"
"Y_GE15","DK0",2012,7.5,"Danmark"
"Y_GE15","DK01",2012,8.2,"Hovedstaden"
"Y_GE15","DK02",2012,6.4,"Sjælland"
"Y_GE15","DK03",2012,7.9,"Syddanmark"
"Y_GE15","DK04",2012,6.8,"Midtjylland"
"Y_GE15","DK05",2012,7.9,"Nordjylland"
"Y_GE15","EA17",2012,11.3,"Euro area (17 countries)"
"Y_GE15","EA18",2012,11.3,"Euro area (18 countries)"
"Y_GE15","EA19",2012,11.4,"Euro area (19 countries)"
"Y_GE15","EE",2012,10,"Estonia"
"Y_GE15","EE0",2012,10,"Eesti"
"Y_GE15","EE00",2012,10,"Eesti"
"Y_GE15","EL",2012,24.4,"Greece"
"Y_GE15","EL3",2012,25.8,"Attiki"
"Y_GE15","EL30",2012,25.8,"Attiki"
"Y_GE15","EL4",2012,20.2,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2012,21.8,"Voreio Aigaio"
"Y_GE15","EL42",2012,15.4,"Notio Aigaio"
"Y_GE15","EL43",2012,22.3,"Kriti"
"Y_GE15","EL5",2012,25.4,"Voreia Ellada"
"Y_GE15","EL51",2012,22.8,"Anatoliki Makedonia, Thraki"
"Y_GE15","EL52",2012,26.2,"Kentriki Makedonia"
"Y_GE15","EL53",2012,29.7,"Dytiki Makedonia"
"Y_GE15","EL54",2012,22.5,"Ipeiros"
"Y_GE15","EL6",2012,23.1,"Kentriki Ellada"
"Y_GE15","EL61",2012,22.6,"Thessalia"
"Y_GE15","EL62",2012,14.7,"Ionia Nisia"
"Y_GE15","EL63",2012,25.6,"Dytiki Ellada"
"Y_GE15","EL64",2012,27.9,"Sterea Ellada"
"Y_GE15","EL65",2012,19.2,"Peloponnisos"
"Y_GE15","ES",2012,24.8,"Spain"
"Y_GE15","ES1",2012,20.5,"Noroeste (ES)"
"Y_GE15","ES11",2012,20.5,"Galicia"
"Y_GE15","ES12",2012,21.8,"Principado de Asturias"
"Y_GE15","ES13",2012,17.8,"Cantabria"
"Y_GE15","ES2",2012,17,"Noreste (ES)"
"Y_GE15","ES21",2012,15.6,"País Vasco"
"Y_GE15","ES22",2012,16.2,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2012,20.6,"La Rioja"
"Y_GE15","ES24",2012,18.7,"Aragón"
"Y_GE15","ES3",2012,18.5,"Comunidad de Madrid"
"Y_GE15","ES30",2012,18.5,"Comunidad de Madrid"
"Y_GE15","ES4",2012,25.6,"Centro (ES)"
"Y_GE15","ES41",2012,19.8,"Castilla y León"
"Y_GE15","ES42",2012,28.6,"Castilla-la Mancha"
"Y_GE15","ES43",2012,33.1,"Extremadura"
"Y_GE15","ES5",2012,24.2,"Este (ES)"
"Y_GE15","ES51",2012,22.5,"Cataluña"
"Y_GE15","ES52",2012,27.2,"Comunidad Valenciana"
"Y_GE15","ES53",2012,23.2,"Illes Balears"
"Y_GE15","ES6",2012,33.3,"Sur (ES)"
"Y_GE15","ES61",2012,34.4,"Andalucía"
"Y_GE15","ES62",2012,27.6,"Región de Murcia"
"Y_GE15","ES63",2012,37,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2012,26.9,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2012,32.6,"Canarias (ES)"
"Y_GE15","ES70",2012,32.6,"Canarias (ES)"
"Y_GE15","EU15",2012,10.6,"European Union (15 countries)"
"Y_GE15","EU27",2012,10.4,"European Union (27 countries)"
"Y_GE15","EU28",2012,10.5,"European Union (28 countries)"
"Y_GE15","FI",2012,7.7,"Finland"
"Y_GE15","FI1",2012,7.7,"Manner-Suomi"
"Y_GE15","FI19",2012,8.2,"Länsi-Suomi"
"Y_GE15","FI1B",2012,6.3,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2012,7.5,"Etelä-Suomi"
"Y_GE15","FI1D",2012,9.5,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2012,NA,"Åland"
"Y_GE15","FI20",2012,NA,"Åland"
"Y_GE15","FR",2012,9.8,"France"
"Y_GE15","FR1",2012,8.1,"Île de France"
"Y_GE15","FR10",2012,8.1,"Île de France"
"Y_GE15","FR2",2012,10.2,"Bassin Parisien"
"Y_GE15","FR21",2012,10.7,"Champagne-Ardenne"
"Y_GE15","FR22",2012,10.6,"Picardie"
"Y_GE15","FR23",2012,10.9,"Haute-Normandie"
"Y_GE15","FR24",2012,10.8,"Centre (FR)"
"Y_GE15","FR25",2012,8.8,"Basse-Normandie"
"Y_GE15","FR26",2012,8.8,"Bourgogne"
"Y_GE15","FR3",2012,13.1,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2012,13.1,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2012,9.9,"Est (FR)"
"Y_GE15","FR41",2012,11.7,"Lorraine"
"Y_GE15","FR42",2012,8.5,"Alsace"
"Y_GE15","FR43",2012,9,"Franche-Comté"
"Y_GE15","FR5",2012,8.2,"Ouest (FR)"
"Y_GE15","FR51",2012,8.4,"Pays de la Loire"
"Y_GE15","FR52",2012,8,"Bretagne"
"Y_GE15","FR53",2012,8.3,"Poitou-Charentes"
"Y_GE15","FR6",2012,8.7,"Sud-Ouest (FR)"
"Y_GE15","FR61",2012,9.4,"Aquitaine"
"Y_GE15","FR62",2012,8.3,"Midi-Pyrénées"
"Y_GE15","FR63",2012,6.7,"Limousin"
"Y_GE15","FR7",2012,8.4,"Centre-Est (FR)"
"Y_GE15","FR71",2012,8,"Rhône-Alpes"
"Y_GE15","FR72",2012,10,"Auvergne"
"Y_GE15","FR8",2012,11.3,"Méditerranée"
"Y_GE15","FR81",2012,15,"Languedoc-Roussillon"
"Y_GE15","FR82",2012,9.6,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2012,7.9,"Corse"
"Y_GE15","FRA",2012,25,"Départements d'outre-mer"
"Y_GE15","FRA1",2012,23,"Guadeloupe"
"Y_GE15","FRA2",2012,21,"Martinique"
"Y_GE15","FRA3",2012,22.3,"Guyane"
"Y_GE15","FRA4",2012,28.6,"La Réunion"
"Y_GE15","HR",2012,15.9,"Croatia"
"Y_GE15","HR0",2012,15.9,"Hrvatska"
"Y_GE15","HR03",2012,14.8,"Jadranska Hrvatska"
"Y_GE15","HR04",2012,16.5,"Kontinentalna Hrvatska"
"Y_GE15","HU",2012,11,"Hungary"
"Y_GE15","HU1",2012,9.5,"Közép-Magyarország"
"Y_GE15","HU10",2012,9.5,"Közép-Magyarország"
"Y_GE15","HU2",2012,9.7,"Dunántúl"
"Y_GE15","HU21",2012,9.9,"Közép-Dunántúl"
"Y_GE15","HU22",2012,7.5,"Nyugat-Dunántúl"
"Y_GE15","HU23",2012,12.1,"Dél-Dunántúl"
"Y_GE15","HU3",2012,13.3,"Alföld és Észak"
"Y_GE15","HU31",2012,16.1,"Észak-Magyarország"
"Y_GE15","HU32",2012,13.9,"Észak-Alföld"
"Y_GE15","HU33",2012,10.3,"Dél-Alföld"
"Y_GE15","IE",2012,14.7,"Ireland"
"Y_GE15","IE0",2012,14.7,"Éire/Ireland"
"Y_GE15","IE01",2012,16.5,"Border, Midland and Western"
"Y_GE15","IE02",2012,14.1,"Southern and Eastern"
"Y_GE15","IS",2012,6,"Iceland"
"Y_GE15","IS0",2012,6,"Ísland"
"Y_GE15","IS00",2012,6,"Ísland"
"Y_GE15","IT",2012,10.7,"Italy"
"Y_GE15","ITC",2012,8,"Nord-Ovest"
"Y_GE15","ITC1",2012,9.2,"Piemonte"
"Y_GE15","ITC2",2012,7.1,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2012,8.1,"Liguria"
"Y_GE15","ITC4",2012,7.4,"Lombardia"
"Y_GE15","ITF",2012,16.9,"Sud"
"Y_GE15","ITF1",2012,10.8,"Abruzzo"
"Y_GE15","ITF2",2012,12,"Molise"
"Y_GE15","ITF3",2012,19.2,"Campania"
"Y_GE15","ITF4",2012,15.7,"Puglia"
"Y_GE15","ITF5",2012,14.5,"Basilicata"
"Y_GE15","ITF6",2012,19.4,"Calabria"
"Y_GE15","ITG",2012,17.5,"Isole"
"Y_GE15","ITG1",2012,18.4,"Sicilia"
"Y_GE15","ITG2",2012,15.4,"Sardegna"
"Y_GE15","ITH",2012,6.6,"Nord-Est"
"Y_GE15","ITH1",2012,4.1,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2012,6.1,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2012,6.4,"Veneto"
"Y_GE15","ITH4",2012,6.7,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2012,7,"Emilia-Romagna"
"Y_GE15","ITI",2012,9.4,"Centro (IT)"
"Y_GE15","ITI1",2012,7.8,"Toscana"
"Y_GE15","ITI2",2012,9.5,"Umbria"
"Y_GE15","ITI3",2012,9.1,"Marche"
"Y_GE15","ITI4",2012,10.6,"Lazio"
"Y_GE15","LT",2012,13.4,"Lithuania"
"Y_GE15","LT0",2012,13.4,"Lietuva"
"Y_GE15","LT00",2012,13.4,"Lietuva"
"Y_GE15","LU",2012,5.1,"Luxembourg"
"Y_GE15","LU0",2012,5.1,"Luxembourg"
"Y_GE15","LU00",2012,5.1,"Luxembourg"
"Y_GE15","LV",2012,15,"Latvia"
"Y_GE15","LV0",2012,15,"Latvija"
"Y_GE15","LV00",2012,15,"Latvija"
"Y_GE15","MK",2012,31,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2012,31,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2012,31,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2012,6.3,"Malta"
"Y_GE15","MT0",2012,6.3,"Malta"
"Y_GE15","MT00",2012,6.3,"Malta"
"Y_GE15","NL",2012,5.8,"Netherlands"
"Y_GE15","NL1",2012,6.6,"Noord-Nederland"
"Y_GE15","NL11",2012,7,"Groningen"
"Y_GE15","NL12",2012,6.4,"Friesland (NL)"
"Y_GE15","NL13",2012,6.4,"Drenthe"
"Y_GE15","NL2",2012,5.6,"Oost-Nederland"
"Y_GE15","NL21",2012,5.6,"Overijssel"
"Y_GE15","NL22",2012,5.3,"Gelderland"
"Y_GE15","NL23",2012,7.3,"Flevoland"
"Y_GE15","NL3",2012,6,"West-Nederland"
"Y_GE15","NL31",2012,5.2,"Utrecht"
"Y_GE15","NL32",2012,5.4,"Noord-Holland"
"Y_GE15","NL33",2012,6.9,"Zuid-Holland"
"Y_GE15","NL34",2012,3.5,"Zeeland"
"Y_GE15","NL4",2012,5.3,"Zuid-Nederland"
"Y_GE15","NL41",2012,5.3,"Noord-Brabant"
"Y_GE15","NL42",2012,5.4,"Limburg (NL)"
"Y_GE15","NO",2012,3.1,"Norway"
"Y_GE15","NO0",2012,3.1,"Norge"
"Y_GE15","NO01",2012,3.2,"Oslo og Akershus"
"Y_GE15","NO02",2012,3,"Hedmark og Oppland"
"Y_GE15","NO03",2012,3.5,"Sør-Østlandet"
"Y_GE15","NO04",2012,2.7,"Agder og Rogaland"
"Y_GE15","NO05",2012,2.9,"Vestlandet"
"Y_GE15","NO06",2012,3.3,"Trøndelag"
"Y_GE15","NO07",2012,3.3,"Nord-Norge"
"Y_GE15","PL",2012,10.1,"Poland"
"Y_GE15","PL1",2012,9,"Region Centralny"
"Y_GE15","PL11",2012,11.1,"Lódzkie"
"Y_GE15","PL12",2012,8,"Mazowieckie"
"Y_GE15","PL2",2012,9.8,"Region Poludniowy"
"Y_GE15","PL21",2012,10.4,"Malopolskie"
"Y_GE15","PL22",2012,9.4,"Slaskie"
"Y_GE15","PL3",2012,11.7,"Region Wschodni"
"Y_GE15","PL31",2012,10.5,"Lubelskie"
"Y_GE15","PL32",2012,13.2,"Podkarpackie"
"Y_GE15","PL33",2012,13.1,"Swietokrzyskie"
"Y_GE15","PL34",2012,9.2,"Podlaskie"
"Y_GE15","PL4",2012,9.2,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2012,8.5,"Wielkopolskie"
"Y_GE15","PL42",2012,10.9,"Zachodniopomorskie"
"Y_GE15","PL43",2012,9,"Lubuskie"
"Y_GE15","PL5",2012,10.7,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2012,11.1,"Dolnoslaskie"
"Y_GE15","PL52",2012,9.5,"Opolskie"
"Y_GE15","PL6",2012,10.7,"Region Pólnocny"
"Y_GE15","PL61",2012,11.9,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2012,11,"Warminsko-Mazurskie"
"Y_GE15","PL63",2012,9.5,"Pomorskie"
"Y_GE15","PT",2012,15.5,"Portugal"
"Y_GE15","PT1",2012,15.5,"Continente"
"Y_GE15","PT11",2012,16,"Norte"
"Y_GE15","PT15",2012,17.6,"Algarve"
"Y_GE15","PT16",2012,11.7,"Centro (PT)"
"Y_GE15","PT17",2012,17.6,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2012,16,"Alentejo"
"Y_GE15","PT2",2012,15.1,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2012,15.1,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2012,17.2,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2012,17.2,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2012,6.8,"Romania"
"Y_GE15","RO1",2012,6.8,"Macroregiunea unu"
"Y_GE15","RO11",2012,4.6,"Nord-Vest"
"Y_GE15","RO12",2012,9.5,"Centru"
"Y_GE15","RO2",2012,6.3,"Macroregiunea doi"
"Y_GE15","RO21",2012,4.2,"Nord-Est"
"Y_GE15","RO22",2012,9.4,"Sud-Est"
"Y_GE15","RO3",2012,8.1,"Macroregiunea trei"
"Y_GE15","RO31",2012,9.5,"Sud - Muntenia"
"Y_GE15","RO32",2012,6.5,"Bucuresti - Ilfov"
"Y_GE15","RO4",2012,5.7,"Macroregiunea patru"
"Y_GE15","RO41",2012,6.1,"Sud-Vest Oltenia"
"Y_GE15","RO42",2012,5.1,"Vest"
"Y_GE15","SE",2012,8,"Sweden"
"Y_GE15","SE1",2012,7.6,"Östra Sverige"
"Y_GE15","SE11",2012,6.8,"Stockholm"
"Y_GE15","SE12",2012,8.6,"Östra Mellansverige"
"Y_GE15","SE2",2012,8.2,"Södra Sverige"
"Y_GE15","SE21",2012,7.4,"Småland med öarna"
"Y_GE15","SE22",2012,9.4,"Sydsverige"
"Y_GE15","SE23",2012,7.7,"Västsverige"
"Y_GE15","SE3",2012,8.3,"Norra Sverige"
"Y_GE15","SE31",2012,8.6,"Norra Mellansverige"
"Y_GE15","SE32",2012,8.4,"Mellersta Norrland"
"Y_GE15","SE33",2012,7.7,"Övre Norrland"
"Y_GE15","SI",2012,8.8,"Slovenia"
"Y_GE15","SI0",2012,8.8,"Slovenija"
"Y_GE15","SI03",2012,9.9,"Vzhodna Slovenija"
"Y_GE15","SI04",2012,7.6,"Zahodna Slovenija"
"Y_GE15","SK",2012,14,"Slovakia"
"Y_GE15","SK0",2012,14,"Slovensko"
"Y_GE15","SK01",2012,5.7,"Bratislavský kraj"
"Y_GE15","SK02",2012,11.3,"Západné Slovensko"
"Y_GE15","SK03",2012,16.2,"Stredné Slovensko"
"Y_GE15","SK04",2012,19,"Východné Slovensko"
"Y_GE15","TR",2012,8.1,"Turkey"
"Y_GE15","TR1",2012,10.7,"Istanbul"
"Y_GE15","TR10",2012,10.7,"Istanbul"
"Y_GE15","TR2",2012,5.4,"Bati Marmara"
"Y_GE15","TR21",2012,6.2,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2012,4.5,"Balikesir, Çanakkale"
"Y_GE15","TR3",2012,8.5,"Ege"
"Y_GE15","TR31",2012,13.3,"Izmir"
"Y_GE15","TR32",2012,6.6,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2012,4.1,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2012,7.6,"Dogu Marmara"
"Y_GE15","TR41",2012,6.4,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2012,8.9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2012,7.3,"Bati Anadolu"
"Y_GE15","TR51",2012,8.3,"Ankara"
"Y_GE15","TR52",2012,5,"Konya, Karaman"
"Y_GE15","TR6",2012,8.5,"Akdeniz"
"Y_GE15","TR61",2012,7.3,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2012,9.1,"Adana, Mersin"
"Y_GE15","TR63",2012,9,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2012,6.9,"Orta Anadolu"
"Y_GE15","TR71",2012,6.2,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2012,7.3,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2012,5.3,"Bati Karadeniz"
"Y_GE15","TR81",2012,6.5,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2012,4.5,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2012,4.9,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2012,5.2,"Dogu Karadeniz"
"Y_GE15","TR90",2012,5.2,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2012,5.9,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2012,5.5,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2012,6.3,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2012,6.6,"Ortadogu Anadolu"
"Y_GE15","TRB1",2012,5.8,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2012,7.5,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2012,11,"Güneydogu Anadolu"
"Y_GE15","TRC1",2012,10.6,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2012,6,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2012,18.8,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2012,7.9,"United Kingdom"
"Y_GE15","UKC",2012,10.1,"North East (UK)"
"Y_GE15","UKC1",2012,11.5,"Tees Valley and Durham"
"Y_GE15","UKC2",2012,9,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2012,8.7,"North West (UK)"
"Y_GE15","UKD1",2012,6.3,"Cumbria"
"Y_GE15","UKD3",2012,10.1,"Greater Manchester"
"Y_GE15","UKD4",2012,7.8,"Lancashire"
"Y_GE15","UKD6",2012,5.9,"Cheshire"
"Y_GE15","UKD7",2012,9.7,"Merseyside"
"Y_GE15","UKE",2012,9,"Yorkshire and The Humber"
"Y_GE15","UKE1",2012,9.7,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2012,5,"North Yorkshire"
"Y_GE15","UKE3",2012,10.4,"South Yorkshire"
"Y_GE15","UKE4",2012,9.4,"West Yorkshire"
"Y_GE15","UKF",2012,7.8,"East Midlands (UK)"
"Y_GE15","UKF1",2012,8.3,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2012,7,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2012,8.5,"Lincolnshire"
"Y_GE15","UKG",2012,8.6,"West Midlands (UK)"
"Y_GE15","UKG1",2012,4.9,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2012,6.7,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2012,11.7,"West Midlands"
"Y_GE15","UKH",2012,6.7,"East of England"
"Y_GE15","UKH1",2012,6.4,"East Anglia"
"Y_GE15","UKH2",2012,6.3,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2012,7.4,"Essex"
"Y_GE15","UKI",2012,9.1,"London"
"Y_GE15","UKI3",2012,6.8,"Inner London - West"
"Y_GE15","UKI4",2012,10.7,"Inner London - East"
"Y_GE15","UKI5",2012,9.5,"Outer London - East and North East"
"Y_GE15","UKI6",2012,7.3,"Outer London - South"
"Y_GE15","UKI7",2012,9.2,"Outer London - West and North West"
"Y_GE15","UKJ",2012,6.3,"South East (UK)"
"Y_GE15","UKJ1",2012,5.7,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2012,5.9,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2012,6.3,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2012,8,"Kent"
"Y_GE15","UKK",2012,5.7,"South West (UK)"
"Y_GE15","UKK1",2012,6.1,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2012,5.1,"Dorset and Somerset"
"Y_GE15","UKK3",2012,5.5,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2012,5.8,"Devon"
"Y_GE15","UKL",2012,8.6,"Wales"
"Y_GE15","UKL1",2012,9.2,"West Wales and The Valleys"
"Y_GE15","UKL2",2012,7.6,"East Wales"
"Y_GE15","UKM",2012,8,"Scotland"
"Y_GE15","UKM2",2012,7.6,"Eastern Scotland"
"Y_GE15","UKM3",2012,9.2,"South Western Scotland"
"Y_GE15","UKM5",2012,4.7,"North Eastern Scotland"
"Y_GE15","UKM6",2012,8.1,"Highlands and Islands"
"Y_GE15","UKN",2012,7.4,"Northern Ireland (UK)"
"Y_GE15","UKN0",2012,7.4,"Northern Ireland (UK)"
"Y_GE25","AT",2012,4.2,"Austria"
"Y_GE25","AT1",2012,5.7,"Ostösterreich"
"Y_GE25","AT11",2012,3.8,"Burgenland (AT)"
"Y_GE25","AT12",2012,4,"Niederösterreich"
"Y_GE25","AT13",2012,7.6,"Wien"
"Y_GE25","AT2",2012,3.7,"Südösterreich"
"Y_GE25","AT21",2012,3.9,"Kärnten"
"Y_GE25","AT22",2012,3.7,"Steiermark"
"Y_GE25","AT3",2012,2.6,"Westösterreich"
"Y_GE25","AT31",2012,2.8,"Oberösterreich"
"Y_GE25","AT32",2012,2.4,"Salzburg"
"Y_GE25","AT33",2012,2.1,"Tirol"
"Y_GE25","AT34",2012,3.1,"Vorarlberg"
"Y_GE25","BE",2012,6.4,"Belgium"
"Y_GE25","BE1",2012,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2012,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2012,3.8,"Vlaams Gewest"
"Y_GE25","BE21",2012,4.7,"Prov. Antwerpen"
"Y_GE25","BE22",2012,3.4,"Prov. Limburg (BE)"
"Y_GE25","BE23",2012,3.4,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2012,3.7,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2012,3.2,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2012,8.3,"Région wallonne"
"Y_GE25","BE31",2012,5.7,"Prov. Brabant Wallon"
"Y_GE25","BE32",2012,10.1,"Prov. Hainaut"
"Y_GE25","BE33",2012,8.9,"Prov. Liège"
"Y_GE25","BE34",2012,5.9,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2012,6,"Prov. Namur"
"Y_GE25","BG",2012,11,"Bulgaria"
"Y_GE25","BG3",2012,12.8,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2012,11,"Severozapaden"
"Y_GE25","BG32",2012,12.9,"Severen tsentralen"
"Y_GE25","BG33",2012,16.6,"Severoiztochen"
"Y_GE25","BG34",2012,10.3,"Yugoiztochen"
"Y_GE25","BG4",2012,9.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2012,7.5,"Yugozapaden"
"Y_GE25","BG42",2012,12.4,"Yuzhen tsentralen"
"Y_GE25","CH",2012,3.5,"Switzerland"
"Y_GE25","CH0",2012,3.5,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2012,5.5,"Région lémanique"
"Y_GE25","CH02",2012,2.8,"Espace Mittelland"
"Y_GE25","CH03",2012,3.4,"Nordwestschweiz"
"Y_GE25","CH04",2012,3.2,"Zürich"
"Y_GE25","CH05",2012,2.9,"Ostschweiz"
"Y_GE25","CH06",2012,2.3,"Zentralschweiz"
"Y_GE25","CH07",2012,5.5,"Ticino"
"Y_GE25","CY",2012,10.1,"Cyprus"
"Y_GE25","CY0",2012,10.1,"Kypros"
"Y_GE25","CY00",2012,10.1,"Kypros"
"Y_GE25","CZ",2012,6,"Czech Republic"
"Y_GE25","CZ0",2012,6,"Ceská republika"
"Y_GE25","CZ01",2012,2.7,"Praha"
"Y_GE25","CZ02",2012,4,"Strední Cechy"
"Y_GE25","CZ03",2012,4.7,"Jihozápad"
"Y_GE25","CZ04",2012,9,"Severozápad"
"Y_GE25","CZ05",2012,6.9,"Severovýchod"
"Y_GE25","CZ06",2012,6.5,"Jihovýchod"
"Y_GE25","CZ07",2012,6.5,"Strední Morava"
"Y_GE25","CZ08",2012,8.6,"Moravskoslezsko"
"Y_GE25","DE",2012,5.1,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2012,3,"Baden-Württemberg"
"Y_GE25","DE11",2012,3.1,"Stuttgart"
"Y_GE25","DE12",2012,3.7,"Karlsruhe"
"Y_GE25","DE13",2012,2.6,"Freiburg"
"Y_GE25","DE14",2012,2.4,"Tübingen"
"Y_GE25","DE2",2012,2.8,"Bayern"
"Y_GE25","DE21",2012,2.5,"Oberbayern"
"Y_GE25","DE22",2012,2.9,"Niederbayern"
"Y_GE25","DE23",2012,2.9,"Oberpfalz"
"Y_GE25","DE24",2012,2.8,"Oberfranken"
"Y_GE25","DE25",2012,3.2,"Mittelfranken"
"Y_GE25","DE26",2012,3.1,"Unterfranken"
"Y_GE25","DE27",2012,2.9,"Schwaben"
"Y_GE25","DE3",2012,10,"Berlin"
"Y_GE25","DE30",2012,10,"Berlin"
"Y_GE25","DE4",2012,7.7,"Brandenburg"
"Y_GE25","DE40",2012,7.7,"Brandenburg"
"Y_GE25","DE5",2012,6,"Bremen"
"Y_GE25","DE50",2012,6,"Bremen"
"Y_GE25","DE6",2012,5.1,"Hamburg"
"Y_GE25","DE60",2012,5.1,"Hamburg"
"Y_GE25","DE7",2012,4.4,"Hessen"
"Y_GE25","DE71",2012,4.4,"Darmstadt"
"Y_GE25","DE72",2012,4.7,"Gießen"
"Y_GE25","DE73",2012,4.1,"Kassel"
"Y_GE25","DE8",2012,10.5,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2012,10.5,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2012,4.5,"Niedersachsen"
"Y_GE25","DE91",2012,5.1,"Braunschweig"
"Y_GE25","DE92",2012,5,"Hannover"
"Y_GE25","DE93",2012,4.1,"Lüneburg"
"Y_GE25","DE94",2012,4,"Weser-Ems"
"Y_GE25","DEA",2012,5.4,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2012,6.1,"Düsseldorf"
"Y_GE25","DEA2",2012,5,"Köln"
"Y_GE25","DEA3",2012,4.5,"Münster"
"Y_GE25","DEA4",2012,4.2,"Detmold"
"Y_GE25","DEA5",2012,6.3,"Arnsberg"
"Y_GE25","DEB",2012,3.6,"Rheinland-Pfalz"
"Y_GE25","DEB1",2012,3.8,"Koblenz"
"Y_GE25","DEB2",2012,2.7,"Trier"
"Y_GE25","DEB3",2012,3.7,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2012,5.5,"Saarland"
"Y_GE25","DEC0",2012,5.5,"Saarland"
"Y_GE25","DED",2012,8.1,"Sachsen"
"Y_GE25","DED2",2012,7.3,"Dresden"
"Y_GE25","DED4",2012,7.8,"Chemnitz"
"Y_GE25","DED5",2012,9.5,"Leipzig"
"Y_GE25","DEE",2012,9.2,"Sachsen-Anhalt"
"Y_GE25","DEE0",2012,9.2,"Sachsen-Anhalt"
"Y_GE25","DEF",2012,4.5,"Schleswig-Holstein"
"Y_GE25","DEF0",2012,4.5,"Schleswig-Holstein"
"Y_GE25","DEG",2012,7.1,"Thüringen"
"Y_GE25","DEG0",2012,7.1,"Thüringen"
"Y_GE25","DK",2012,6.3,"Denmark"
"Y_GE25","DK0",2012,6.3,"Danmark"
"Y_GE25","DK01",2012,7.1,"Hovedstaden"
"Y_GE25","DK02",2012,5,"Sjælland"
"Y_GE25","DK03",2012,6.6,"Syddanmark"
"Y_GE25","DK04",2012,5.6,"Midtjylland"
"Y_GE25","DK05",2012,6.7,"Nordjylland"
"Y_GE25","EA17",2012,10,"Euro area (17 countries)"
"Y_GE25","EA18",2012,10.1,"Euro area (18 countries)"
"Y_GE25","EA19",2012,10.1,"Euro area (19 countries)"
"Y_GE25","EE",2012,8.9,"Estonia"
"Y_GE25","EE0",2012,8.9,"Eesti"
"Y_GE25","EE00",2012,8.9,"Eesti"
"Y_GE25","EL",2012,22.2,"Greece"
"Y_GE25","EL3",2012,23.7,"Attiki"
"Y_GE25","EL30",2012,23.7,"Attiki"
"Y_GE25","EL4",2012,18.3,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2012,19.4,"Voreio Aigaio"
"Y_GE25","EL42",2012,13.5,"Notio Aigaio"
"Y_GE25","EL43",2012,20.5,"Kriti"
"Y_GE25","EL5",2012,23,"Voreia Ellada"
"Y_GE25","EL51",2012,20.2,"Anatoliki Makedonia, Thraki"
"Y_GE25","EL52",2012,24.1,"Kentriki Makedonia"
"Y_GE25","EL53",2012,26.4,"Dytiki Makedonia"
"Y_GE25","EL54",2012,19.5,"Ipeiros"
"Y_GE25","EL6",2012,20.7,"Kentriki Ellada"
"Y_GE25","EL61",2012,20.3,"Thessalia"
"Y_GE25","EL62",2012,14.2,"Ionia Nisia"
"Y_GE25","EL63",2012,23.2,"Dytiki Ellada"
"Y_GE25","EL64",2012,25.1,"Sterea Ellada"
"Y_GE25","EL65",2012,16.7,"Peloponnisos"
"Y_GE25","ES",2012,22.4,"Spain"
"Y_GE25","ES1",2012,18.9,"Noroeste (ES)"
"Y_GE25","ES11",2012,18.9,"Galicia"
"Y_GE25","ES12",2012,20.4,"Principado de Asturias"
"Y_GE25","ES13",2012,16.5,"Cantabria"
"Y_GE25","ES2",2012,15.2,"Noreste (ES)"
"Y_GE25","ES21",2012,14,"País Vasco"
"Y_GE25","ES22",2012,14.5,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2012,18.3,"La Rioja"
"Y_GE25","ES24",2012,16.9,"Aragón"
"Y_GE25","ES3",2012,16.4,"Comunidad de Madrid"
"Y_GE25","ES30",2012,16.4,"Comunidad de Madrid"
"Y_GE25","ES4",2012,23.1,"Centro (ES)"
"Y_GE25","ES41",2012,17.8,"Castilla y León"
"Y_GE25","ES42",2012,26,"Castilla-la Mancha"
"Y_GE25","ES43",2012,29.9,"Extremadura"
"Y_GE25","ES5",2012,21.9,"Este (ES)"
"Y_GE25","ES51",2012,20.1,"Cataluña"
"Y_GE25","ES52",2012,25,"Comunidad Valenciana"
"Y_GE25","ES53",2012,20.8,"Illes Balears"
"Y_GE25","ES6",2012,30.6,"Sur (ES)"
"Y_GE25","ES61",2012,31.6,"Andalucía"
"Y_GE25","ES62",2012,25.4,"Región de Murcia"
"Y_GE25","ES63",2012,33.4,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2012,23.7,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2012,29.9,"Canarias (ES)"
"Y_GE25","ES70",2012,29.9,"Canarias (ES)"
"Y_GE25","EU15",2012,9.2,"European Union (15 countries)"
"Y_GE25","EU27",2012,9,"European Union (27 countries)"
"Y_GE25","EU28",2012,9,"European Union (28 countries)"
"Y_GE25","FI",2012,6.1,"Finland"
"Y_GE25","FI1",2012,6.1,"Manner-Suomi"
"Y_GE25","FI19",2012,6.2,"Länsi-Suomi"
"Y_GE25","FI1B",2012,5,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2012,6.1,"Etelä-Suomi"
"Y_GE25","FI1D",2012,7.7,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2012,NA,"Åland"
"Y_GE25","FI20",2012,NA,"Åland"
"Y_GE25","FR",2012,8.2,"France"
"Y_GE25","FR1",2012,7.1,"Île de France"
"Y_GE25","FR10",2012,7.1,"Île de France"
"Y_GE25","FR2",2012,8.3,"Bassin Parisien"
"Y_GE25","FR21",2012,8.9,"Champagne-Ardenne"
"Y_GE25","FR22",2012,8.8,"Picardie"
"Y_GE25","FR23",2012,8.9,"Haute-Normandie"
"Y_GE25","FR24",2012,8.6,"Centre (FR)"
"Y_GE25","FR25",2012,7.2,"Basse-Normandie"
"Y_GE25","FR26",2012,7.1,"Bourgogne"
"Y_GE25","FR3",2012,10.3,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2012,10.3,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2012,8.3,"Est (FR)"
"Y_GE25","FR41",2012,10,"Lorraine"
"Y_GE25","FR42",2012,6.8,"Alsace"
"Y_GE25","FR43",2012,7.7,"Franche-Comté"
"Y_GE25","FR5",2012,6.8,"Ouest (FR)"
"Y_GE25","FR51",2012,6.7,"Pays de la Loire"
"Y_GE25","FR52",2012,7.1,"Bretagne"
"Y_GE25","FR53",2012,6.6,"Poitou-Charentes"
"Y_GE25","FR6",2012,7.5,"Sud-Ouest (FR)"
"Y_GE25","FR61",2012,8,"Aquitaine"
"Y_GE25","FR62",2012,7.5,"Midi-Pyrénées"
"Y_GE25","FR63",2012,5.7,"Limousin"
"Y_GE25","FR7",2012,6.9,"Centre-Est (FR)"
"Y_GE25","FR71",2012,6.7,"Rhône-Alpes"
"Y_GE25","FR72",2012,7.8,"Auvergne"
"Y_GE25","FR8",2012,9.6,"Méditerranée"
"Y_GE25","FR81",2012,12.3,"Languedoc-Roussillon"
"Y_GE25","FR82",2012,8.4,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2012,NA,"Corse"
"Y_GE25","FRA",2012,21.7,"Départements d'outre-mer"
"Y_GE25","FRA1",2012,20.6,"Guadeloupe"
"Y_GE25","FRA2",2012,18.1,"Martinique"
"Y_GE25","FRA3",2012,18.9,"Guyane"
"Y_GE25","FRA4",2012,24.7,"La Réunion"
"Y_GE25","HR",2012,13.6,"Croatia"
"Y_GE25","HR0",2012,13.6,"Hrvatska"
"Y_GE25","HR03",2012,12.9,"Jadranska Hrvatska"
"Y_GE25","HR04",2012,14,"Kontinentalna Hrvatska"
"Y_GE25","HU",2012,9.7,"Hungary"
"Y_GE25","HU1",2012,8.6,"Közép-Magyarország"
"Y_GE25","HU10",2012,8.6,"Közép-Magyarország"
"Y_GE25","HU2",2012,8.5,"Dunántúl"
"Y_GE25","HU21",2012,8.7,"Közép-Dunántúl"
"Y_GE25","HU22",2012,6.4,"Nyugat-Dunántúl"
"Y_GE25","HU23",2012,10.8,"Dél-Dunántúl"
"Y_GE25","HU3",2012,11.6,"Alföld és Észak"
"Y_GE25","HU31",2012,14.1,"Észak-Magyarország"
"Y_GE25","HU32",2012,12,"Észak-Alföld"
"Y_GE25","HU33",2012,8.9,"Dél-Alföld"
"Y_GE25","IE",2012,12.8,"Ireland"
"Y_GE25","IE0",2012,12.8,"Éire/Ireland"
"Y_GE25","IE01",2012,14.4,"Border, Midland and Western"
"Y_GE25","IE02",2012,12.3,"Southern and Eastern"
"Y_GE25","IS",2012,4.4,"Iceland"
"Y_GE25","IS0",2012,4.4,"Ísland"
"Y_GE25","IS00",2012,4.4,"Ísland"
"Y_GE25","IT",2012,8.9,"Italy"
"Y_GE25","ITC",2012,6.6,"Nord-Ovest"
"Y_GE25","ITC1",2012,7.6,"Piemonte"
"Y_GE25","ITC2",2012,5.8,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2012,6.7,"Liguria"
"Y_GE25","ITC4",2012,6.1,"Lombardia"
"Y_GE25","ITF",2012,14.3,"Sud"
"Y_GE25","ITF1",2012,9,"Abruzzo"
"Y_GE25","ITF2",2012,9.9,"Molise"
"Y_GE25","ITF3",2012,16.5,"Campania"
"Y_GE25","ITF4",2012,13.3,"Puglia"
"Y_GE25","ITF5",2012,11.8,"Basilicata"
"Y_GE25","ITF6",2012,16.4,"Calabria"
"Y_GE25","ITG",2012,14.6,"Isole"
"Y_GE25","ITG1",2012,15.3,"Sicilia"
"Y_GE25","ITG2",2012,13,"Sardegna"
"Y_GE25","ITH",2012,5.4,"Nord-Est"
"Y_GE25","ITH1",2012,3.3,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2012,5,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2012,5.2,"Veneto"
"Y_GE25","ITH4",2012,5.5,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2012,5.8,"Emilia-Romagna"
"Y_GE25","ITI",2012,7.8,"Centro (IT)"
"Y_GE25","ITI1",2012,6.5,"Toscana"
"Y_GE25","ITI2",2012,7.7,"Umbria"
"Y_GE25","ITI3",2012,7.8,"Marche"
"Y_GE25","ITI4",2012,8.8,"Lazio"
"Y_GE25","LT",2012,12.2,"Lithuania"
"Y_GE25","LT0",2012,12.2,"Lietuva"
"Y_GE25","LT00",2012,12.2,"Lietuva"
"Y_GE25","LU",2012,4.2,"Luxembourg"
"Y_GE25","LU0",2012,4.2,"Luxembourg"
"Y_GE25","LU00",2012,4.2,"Luxembourg"
"Y_GE25","LV",2012,13.6,"Latvia"
"Y_GE25","LV0",2012,13.6,"Latvija"
"Y_GE25","LV00",2012,13.6,"Latvija"
"Y_GE25","MK",2012,28.2,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2012,28.2,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2012,28.2,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2012,4.9,"Malta"
"Y_GE25","MT0",2012,4.9,"Malta"
"Y_GE25","MT00",2012,4.9,"Malta"
"Y_GE25","NL",2012,4.7,"Netherlands"
"Y_GE25","NL1",2012,5.3,"Noord-Nederland"
"Y_GE25","NL11",2012,5.3,"Groningen"
"Y_GE25","NL12",2012,5.3,"Friesland (NL)"
"Y_GE25","NL13",2012,5.3,"Drenthe"
"Y_GE25","NL2",2012,4.5,"Oost-Nederland"
"Y_GE25","NL21",2012,4.5,"Overijssel"
"Y_GE25","NL22",2012,4.3,"Gelderland"
"Y_GE25","NL23",2012,5.9,"Flevoland"
"Y_GE25","NL3",2012,4.9,"West-Nederland"
"Y_GE25","NL31",2012,4.1,"Utrecht"
"Y_GE25","NL32",2012,4.5,"Noord-Holland"
"Y_GE25","NL33",2012,5.6,"Zuid-Holland"
"Y_GE25","NL34",2012,2.8,"Zeeland"
"Y_GE25","NL4",2012,4.3,"Zuid-Nederland"
"Y_GE25","NL41",2012,4.2,"Noord-Brabant"
"Y_GE25","NL42",2012,4.4,"Limburg (NL)"
"Y_GE25","NO",2012,2.3,"Norway"
"Y_GE25","NO0",2012,2.3,"Norge"
"Y_GE25","NO01",2012,2.4,"Oslo og Akershus"
"Y_GE25","NO02",2012,2.5,"Hedmark og Oppland"
"Y_GE25","NO03",2012,2.5,"Sør-Østlandet"
"Y_GE25","NO04",2012,2,"Agder og Rogaland"
"Y_GE25","NO05",2012,1.9,"Vestlandet"
"Y_GE25","NO06",2012,2.4,"Trøndelag"
"Y_GE25","NO07",2012,2.2,"Nord-Norge"
"Y_GE25","PL",2012,8.5,"Poland"
"Y_GE25","PL1",2012,7.8,"Region Centralny"
"Y_GE25","PL11",2012,9.6,"Lódzkie"
"Y_GE25","PL12",2012,7,"Mazowieckie"
"Y_GE25","PL2",2012,8.3,"Region Poludniowy"
"Y_GE25","PL21",2012,8.4,"Malopolskie"
"Y_GE25","PL22",2012,8.2,"Slaskie"
"Y_GE25","PL3",2012,9.6,"Region Wschodni"
"Y_GE25","PL31",2012,8.6,"Lubelskie"
"Y_GE25","PL32",2012,10.6,"Podkarpackie"
"Y_GE25","PL33",2012,11.2,"Swietokrzyskie"
"Y_GE25","PL34",2012,7.8,"Podlaskie"
"Y_GE25","PL4",2012,7.5,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2012,6.8,"Wielkopolskie"
"Y_GE25","PL42",2012,9.1,"Zachodniopomorskie"
"Y_GE25","PL43",2012,7.4,"Lubuskie"
"Y_GE25","PL5",2012,9,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2012,9.3,"Dolnoslaskie"
"Y_GE25","PL52",2012,8.1,"Opolskie"
"Y_GE25","PL6",2012,9,"Region Pólnocny"
"Y_GE25","PL61",2012,9.8,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2012,9.4,"Warminsko-Mazurskie"
"Y_GE25","PL63",2012,8,"Pomorskie"
"Y_GE25","PT",2012,13.6,"Portugal"
"Y_GE25","PT1",2012,13.7,"Continente"
"Y_GE25","PT11",2012,14.4,"Norte"
"Y_GE25","PT15",2012,15.9,"Algarve"
"Y_GE25","PT16",2012,9.9,"Centro (PT)"
"Y_GE25","PT17",2012,15.5,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2012,13.8,"Alentejo"
"Y_GE25","PT2",2012,12.1,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2012,12.1,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2012,14.3,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2012,14.3,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2012,5.4,"Romania"
"Y_GE25","RO1",2012,5.3,"Macroregiunea unu"
"Y_GE25","RO11",2012,3.6,"Nord-Vest"
"Y_GE25","RO12",2012,7.5,"Centru"
"Y_GE25","RO2",2012,5.1,"Macroregiunea doi"
"Y_GE25","RO21",2012,3.4,"Nord-Est"
"Y_GE25","RO22",2012,7.6,"Sud-Est"
"Y_GE25","RO3",2012,6.5,"Macroregiunea trei"
"Y_GE25","RO31",2012,7.5,"Sud - Muntenia"
"Y_GE25","RO32",2012,5.3,"Bucuresti - Ilfov"
"Y_GE25","RO4",2012,4.5,"Macroregiunea patru"
"Y_GE25","RO41",2012,5,"Sud-Vest Oltenia"
"Y_GE25","RO42",2012,3.7,"Vest"
"Y_GE25","SE",2012,5.7,"Sweden"
"Y_GE25","SE1",2012,5.4,"Östra Sverige"
"Y_GE25","SE11",2012,4.9,"Stockholm"
"Y_GE25","SE12",2012,6.1,"Östra Mellansverige"
"Y_GE25","SE2",2012,5.9,"Södra Sverige"
"Y_GE25","SE21",2012,5.1,"Småland med öarna"
"Y_GE25","SE22",2012,7,"Sydsverige"
"Y_GE25","SE23",2012,5.4,"Västsverige"
"Y_GE25","SE3",2012,5.7,"Norra Sverige"
"Y_GE25","SE31",2012,6.2,"Norra Mellansverige"
"Y_GE25","SE32",2012,5.7,"Mellersta Norrland"
"Y_GE25","SE33",2012,5.1,"Övre Norrland"
"Y_GE25","SI",2012,7.9,"Slovenia"
"Y_GE25","SI0",2012,7.9,"Slovenija"
"Y_GE25","SI03",2012,8.9,"Vzhodna Slovenija"
"Y_GE25","SI04",2012,6.7,"Zahodna Slovenija"
"Y_GE25","SK",2012,12.2,"Slovakia"
"Y_GE25","SK0",2012,12.2,"Slovensko"
"Y_GE25","SK01",2012,5,"Bratislavský kraj"
"Y_GE25","SK02",2012,10.2,"Západné Slovensko"
"Y_GE25","SK03",2012,13.9,"Stredné Slovensko"
"Y_GE25","SK04",2012,16.5,"Východné Slovensko"
"Y_GE25","TR",2012,6.7,"Turkey"
"Y_GE25","TR1",2012,9,"Istanbul"
"Y_GE25","TR10",2012,9,"Istanbul"
"Y_GE25","TR2",2012,4.1,"Bati Marmara"
"Y_GE25","TR21",2012,4.8,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2012,3.4,"Balikesir, Çanakkale"
"Y_GE25","TR3",2012,7.2,"Ege"
"Y_GE25","TR31",2012,11.4,"Izmir"
"Y_GE25","TR32",2012,5.5,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2012,3.2,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2012,6.2,"Dogu Marmara"
"Y_GE25","TR41",2012,5.3,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2012,7.2,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2012,5.7,"Bati Anadolu"
"Y_GE25","TR51",2012,6.5,"Ankara"
"Y_GE25","TR52",2012,3.8,"Konya, Karaman"
"Y_GE25","TR6",2012,7.2,"Akdeniz"
"Y_GE25","TR61",2012,6.3,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2012,7.7,"Adana, Mersin"
"Y_GE25","TR63",2012,7.5,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2012,5.6,"Orta Anadolu"
"Y_GE25","TR71",2012,4.4,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2012,6.3,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2012,4.4,"Bati Karadeniz"
"Y_GE25","TR81",2012,5.1,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2012,3.8,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2012,4.3,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2012,3.6,"Dogu Karadeniz"
"Y_GE25","TR90",2012,3.6,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2012,4.9,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2012,4.6,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2012,5.2,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2012,5.2,"Ortadogu Anadolu"
"Y_GE25","TRB1",2012,4.3,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2012,6.2,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2012,9.5,"Güneydogu Anadolu"
"Y_GE25","TRC1",2012,9.6,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2012,5.5,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2012,15.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2012,5.7,"United Kingdom"
"Y_GE25","UKC",2012,7.4,"North East (UK)"
"Y_GE25","UKC1",2012,8,"Tees Valley and Durham"
"Y_GE25","UKC2",2012,6.9,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2012,6,"North West (UK)"
"Y_GE25","UKD1",2012,5,"Cumbria"
"Y_GE25","UKD3",2012,7.2,"Greater Manchester"
"Y_GE25","UKD4",2012,4.8,"Lancashire"
"Y_GE25","UKD6",2012,4.2,"Cheshire"
"Y_GE25","UKD7",2012,6.7,"Merseyside"
"Y_GE25","UKE",2012,6.4,"Yorkshire and The Humber"
"Y_GE25","UKE1",2012,7.3,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2012,3.1,"North Yorkshire"
"Y_GE25","UKE3",2012,8,"South Yorkshire"
"Y_GE25","UKE4",2012,6.4,"West Yorkshire"
"Y_GE25","UKF",2012,5.6,"East Midlands (UK)"
"Y_GE25","UKF1",2012,5.8,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2012,5.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2012,6.3,"Lincolnshire"
"Y_GE25","UKG",2012,6.1,"West Midlands (UK)"
"Y_GE25","UKG1",2012,3.2,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2012,4.5,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2012,8.6,"West Midlands"
"Y_GE25","UKH",2012,4.9,"East of England"
"Y_GE25","UKH1",2012,4.6,"East Anglia"
"Y_GE25","UKH2",2012,5.2,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2012,5.1,"Essex"
"Y_GE25","UKI",2012,7,"London"
"Y_GE25","UKI3",2012,5.5,"Inner London - West"
"Y_GE25","UKI4",2012,8.2,"Inner London - East"
"Y_GE25","UKI5",2012,7.2,"Outer London - East and North East"
"Y_GE25","UKI6",2012,5.5,"Outer London - South"
"Y_GE25","UKI7",2012,7.3,"Outer London - West and North West"
"Y_GE25","UKJ",2012,4.5,"South East (UK)"
"Y_GE25","UKJ1",2012,4.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2012,4,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2012,4.7,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2012,5.3,"Kent"
"Y_GE25","UKK",2012,4,"South West (UK)"
"Y_GE25","UKK1",2012,4.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2012,3.9,"Dorset and Somerset"
"Y_GE25","UKK3",2012,4.1,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2012,3.6,"Devon"
"Y_GE25","UKL",2012,5.8,"Wales"
"Y_GE25","UKL1",2012,6.7,"West Wales and The Valleys"
"Y_GE25","UKL2",2012,4.4,"East Wales"
"Y_GE25","UKM",2012,5.4,"Scotland"
"Y_GE25","UKM2",2012,5,"Eastern Scotland"
"Y_GE25","UKM3",2012,6.2,"South Western Scotland"
"Y_GE25","UKM5",2012,3.3,"North Eastern Scotland"
"Y_GE25","UKM6",2012,6,"Highlands and Islands"
"Y_GE25","UKN",2012,5.7,"Northern Ireland (UK)"
"Y_GE25","UKN0",2012,5.7,"Northern Ireland (UK)"
"Y15-24","AT",2011,8.9,"Austria"
"Y15-24","AT1",2011,12.8,"Ostösterreich"
"Y15-24","AT11",2011,NA,"Burgenland (AT)"
"Y15-24","AT12",2011,9.4,"Niederösterreich"
"Y15-24","AT13",2011,17.3,"Wien"
"Y15-24","AT2",2011,6.3,"Südösterreich"
"Y15-24","AT21",2011,8.7,"Kärnten"
"Y15-24","AT22",2011,5.3,"Steiermark"
"Y15-24","AT3",2011,6.8,"Westösterreich"
"Y15-24","AT31",2011,7.1,"Oberösterreich"
"Y15-24","AT32",2011,NA,"Salzburg"
"Y15-24","AT33",2011,NA,"Tirol"
"Y15-24","AT34",2011,NA,"Vorarlberg"
"Y15-24","BE",2011,18.7,"Belgium"
"Y15-24","BE1",2011,35.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2011,35.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2011,12.7,"Vlaams Gewest"
"Y15-24","BE21",2011,15.8,"Prov. Antwerpen"
"Y15-24","BE22",2011,12.6,"Prov. Limburg (BE)"
"Y15-24","BE23",2011,11.4,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2011,10.4,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2011,11.4,"Prov. West-Vlaanderen"
"Y15-24","BE3",2011,25.2,"Région wallonne"
"Y15-24","BE31",2011,22.3,"Prov. Brabant Wallon"
"Y15-24","BE32",2011,30.8,"Prov. Hainaut"
"Y15-24","BE33",2011,22.5,"Prov. Liège"
"Y15-24","BE34",2011,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2011,22,"Prov. Namur"
"Y15-24","BG",2011,25,"Bulgaria"
"Y15-24","BG3",2011,29.7,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2011,31.8,"Severozapaden"
"Y15-24","BG32",2011,29.4,"Severen tsentralen"
"Y15-24","BG33",2011,30.1,"Severoiztochen"
"Y15-24","BG34",2011,28,"Yugoiztochen"
"Y15-24","BG4",2011,20.9,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2011,16,"Yugozapaden"
"Y15-24","BG42",2011,31.6,"Yuzhen tsentralen"
"Y15-24","CH",2011,7.7,"Switzerland"
"Y15-24","CH0",2011,7.7,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2011,13.2,"Région lémanique"
"Y15-24","CH02",2011,7.1,"Espace Mittelland"
"Y15-24","CH03",2011,7.1,"Nordwestschweiz"
"Y15-24","CH04",2011,4.3,"Zürich"
"Y15-24","CH05",2011,6.8,"Ostschweiz"
"Y15-24","CH06",2011,4.2,"Zentralschweiz"
"Y15-24","CH07",2011,17.3,"Ticino"
"Y15-24","CY",2011,22.4,"Cyprus"
"Y15-24","CY0",2011,22.4,"Kypros"
"Y15-24","CY00",2011,22.4,"Kypros"
"Y15-24","CZ",2011,18.1,"Czech Republic"
"Y15-24","CZ0",2011,18.1,"Ceská republika"
"Y15-24","CZ01",2011,10.1,"Praha"
"Y15-24","CZ02",2011,16.1,"Strední Cechy"
"Y15-24","CZ03",2011,14.2,"Jihozápad"
"Y15-24","CZ04",2011,26.9,"Severozápad"
"Y15-24","CZ05",2011,17.9,"Severovýchod"
"Y15-24","CZ06",2011,18.9,"Jihovýchod"
"Y15-24","CZ07",2011,20.2,"Strední Morava"
"Y15-24","CZ08",2011,18.3,"Moravskoslezsko"
"Y15-24","DE",2011,8.5,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2011,5.6,"Baden-Württemberg"
"Y15-24","DE11",2011,6.2,"Stuttgart"
"Y15-24","DE12",2011,6.6,"Karlsruhe"
"Y15-24","DE13",2011,4.8,"Freiburg"
"Y15-24","DE14",2011,NA,"Tübingen"
"Y15-24","DE2",2011,5.4,"Bayern"
"Y15-24","DE21",2011,4.5,"Oberbayern"
"Y15-24","DE22",2011,NA,"Niederbayern"
"Y15-24","DE23",2011,NA,"Oberpfalz"
"Y15-24","DE24",2011,NA,"Oberfranken"
"Y15-24","DE25",2011,6.3,"Mittelfranken"
"Y15-24","DE26",2011,NA,"Unterfranken"
"Y15-24","DE27",2011,6.7,"Schwaben"
"Y15-24","DE3",2011,13.3,"Berlin"
"Y15-24","DE30",2011,13.3,"Berlin"
"Y15-24","DE4",2011,12.4,"Brandenburg"
"Y15-24","DE40",2011,12.4,"Brandenburg"
"Y15-24","DE5",2011,15.3,"Bremen"
"Y15-24","DE50",2011,15.3,"Bremen"
"Y15-24","DE6",2011,6.6,"Hamburg"
"Y15-24","DE60",2011,6.6,"Hamburg"
"Y15-24","DE7",2011,8.5,"Hessen"
"Y15-24","DE71",2011,9,"Darmstadt"
"Y15-24","DE72",2011,9.6,"Gießen"
"Y15-24","DE73",2011,NA,"Kassel"
"Y15-24","DE8",2011,10.7,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2011,10.7,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2011,9.5,"Niedersachsen"
"Y15-24","DE91",2011,11,"Braunschweig"
"Y15-24","DE92",2011,11.9,"Hannover"
"Y15-24","DE93",2011,9.3,"Lüneburg"
"Y15-24","DE94",2011,6.7,"Weser-Ems"
"Y15-24","DEA",2011,9.7,"Nordrhein-Westfalen"
"Y15-24","DEA1",2011,11.7,"Düsseldorf"
"Y15-24","DEA2",2011,9.5,"Köln"
"Y15-24","DEA3",2011,7,"Münster"
"Y15-24","DEA4",2011,9.1,"Detmold"
"Y15-24","DEA5",2011,9.6,"Arnsberg"
"Y15-24","DEB",2011,9.3,"Rheinland-Pfalz"
"Y15-24","DEB1",2011,7.6,"Koblenz"
"Y15-24","DEB2",2011,NA,"Trier"
"Y15-24","DEB3",2011,10.6,"Rheinhessen-Pfalz"
"Y15-24","DEC",2011,10.3,"Saarland"
"Y15-24","DEC0",2011,10.3,"Saarland"
"Y15-24","DED",2011,10.3,"Sachsen"
"Y15-24","DED2",2011,9.8,"Dresden"
"Y15-24","DED4",2011,9.6,"Chemnitz"
"Y15-24","DED5",2011,11.8,"Leipzig"
"Y15-24","DEE",2011,14,"Sachsen-Anhalt"
"Y15-24","DEE0",2011,14,"Sachsen-Anhalt"
"Y15-24","DEF",2011,9,"Schleswig-Holstein"
"Y15-24","DEF0",2011,9,"Schleswig-Holstein"
"Y15-24","DEG",2011,8.2,"Thüringen"
"Y15-24","DEG0",2011,8.2,"Thüringen"
"Y15-24","DK",2011,14.2,"Denmark"
"Y15-24","DK0",2011,14.2,"Danmark"
"Y15-24","DK01",2011,15.4,"Hovedstaden"
"Y15-24","DK02",2011,15,"Sjælland"
"Y15-24","DK03",2011,14.2,"Syddanmark"
"Y15-24","DK04",2011,12.5,"Midtjylland"
"Y15-24","DK05",2011,13.9,"Nordjylland"
"Y15-24","EA17",2011,21.2,"Euro area (17 countries)"
"Y15-24","EA18",2011,21.3,"Euro area (18 countries)"
"Y15-24","EA19",2011,21.4,"Euro area (19 countries)"
"Y15-24","EE",2011,22.4,"Estonia"
"Y15-24","EE0",2011,22.4,"Eesti"
"Y15-24","EE00",2011,22.4,"Eesti"
"Y15-24","EL",2011,44.7,"Greece"
"Y15-24","EL3",2011,43.2,"Attiki"
"Y15-24","EL30",2011,43.2,"Attiki"
"Y15-24","EL4",2011,39.3,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2011,43,"Voreio Aigaio"
"Y15-24","EL42",2011,36.8,"Notio Aigaio"
"Y15-24","EL43",2011,39.8,"Kriti"
"Y15-24","EL5",2011,51.3,"Voreia Ellada"
"Y15-24","EL51",2011,51.8,"Anatoliki Makedonia, Thraki"
"Y15-24","EL52",2011,51.4,"Kentriki Makedonia"
"Y15-24","EL53",2011,52.7,"Dytiki Makedonia"
"Y15-24","EL54",2011,48.6,"Ipeiros"
"Y15-24","EL6",2011,42.9,"Kentriki Ellada"
"Y15-24","EL61",2011,46.7,"Thessalia"
"Y15-24","EL62",2011,26.2,"Ionia Nisia"
"Y15-24","EL63",2011,45.1,"Dytiki Ellada"
"Y15-24","EL64",2011,42.5,"Sterea Ellada"
"Y15-24","EL65",2011,39,"Peloponnisos"
"Y15-24","ES",2011,46.2,"Spain"
"Y15-24","ES1",2011,40.3,"Noroeste (ES)"
"Y15-24","ES11",2011,37.7,"Galicia"
"Y15-24","ES12",2011,48.5,"Principado de Asturias"
"Y15-24","ES13",2011,40.6,"Cantabria"
"Y15-24","ES2",2011,36.2,"Noreste (ES)"
"Y15-24","ES21",2011,34.1,"País Vasco"
"Y15-24","ES22",2011,29.3,"Comunidad Foral de Navarra"
"Y15-24","ES23",2011,46.1,"La Rioja"
"Y15-24","ES24",2011,39.9,"Aragón"
"Y15-24","ES3",2011,40.8,"Comunidad de Madrid"
"Y15-24","ES30",2011,40.8,"Comunidad de Madrid"
"Y15-24","ES4",2011,45,"Centro (ES)"
"Y15-24","ES41",2011,38.6,"Castilla y León"
"Y15-24","ES42",2011,47.7,"Castilla-la Mancha"
"Y15-24","ES43",2011,51,"Extremadura"
"Y15-24","ES5",2011,46.4,"Este (ES)"
"Y15-24","ES51",2011,43.8,"Cataluña"
"Y15-24","ES52",2011,51.4,"Comunidad Valenciana"
"Y15-24","ES53",2011,42.7,"Illes Balears"
"Y15-24","ES6",2011,53.3,"Sur (ES)"
"Y15-24","ES61",2011,54.1,"Andalucía"
"Y15-24","ES62",2011,48,"Región de Murcia"
"Y15-24","ES63",2011,63.9,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2011,63.8,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2011,50.8,"Canarias (ES)"
"Y15-24","ES70",2011,50.8,"Canarias (ES)"
"Y15-24","EU15",2011,21,"European Union (15 countries)"
"Y15-24","EU27",2011,21.7,"European Union (27 countries)"
"Y15-24","EU28",2011,21.8,"European Union (28 countries)"
"Y15-24","FI",2011,20.1,"Finland"
"Y15-24","FI1",2011,20.1,"Manner-Suomi"
"Y15-24","FI19",2011,23.1,"Länsi-Suomi"
"Y15-24","FI1B",2011,14.5,"Helsinki-Uusimaa"
"Y15-24","FI1C",2011,21.5,"Etelä-Suomi"
"Y15-24","FI1D",2011,23.3,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2011,NA,"Åland"
"Y15-24","FI20",2011,NA,"Åland"
"Y15-24","FR",2011,22.9,"France"
"Y15-24","FR1",2011,19.1,"Île de France"
"Y15-24","FR10",2011,19.1,"Île de France"
"Y15-24","FR2",2011,22.9,"Bassin Parisien"
"Y15-24","FR21",2011,26.6,"Champagne-Ardenne"
"Y15-24","FR22",2011,23.5,"Picardie"
"Y15-24","FR23",2011,22,"Haute-Normandie"
"Y15-24","FR24",2011,20.2,"Centre (FR)"
"Y15-24","FR25",2011,24,"Basse-Normandie"
"Y15-24","FR26",2011,23.3,"Bourgogne"
"Y15-24","FR3",2011,30.6,"Nord - Pas-de-Calais"
"Y15-24","FR30",2011,30.6,"Nord - Pas-de-Calais"
"Y15-24","FR4",2011,20.7,"Est (FR)"
"Y15-24","FR41",2011,21,"Lorraine"
"Y15-24","FR42",2011,21.4,"Alsace"
"Y15-24","FR43",2011,18.5,"Franche-Comté"
"Y15-24","FR5",2011,18.7,"Ouest (FR)"
"Y15-24","FR51",2011,17.6,"Pays de la Loire"
"Y15-24","FR52",2011,18.8,"Bretagne"
"Y15-24","FR53",2011,21.3,"Poitou-Charentes"
"Y15-24","FR6",2011,22.9,"Sud-Ouest (FR)"
"Y15-24","FR61",2011,24.9,"Aquitaine"
"Y15-24","FR62",2011,21.3,"Midi-Pyrénées"
"Y15-24","FR63",2011,21.2,"Limousin"
"Y15-24","FR7",2011,20.2,"Centre-Est (FR)"
"Y15-24","FR71",2011,19.6,"Rhône-Alpes"
"Y15-24","FR72",2011,23.3,"Auvergne"
"Y15-24","FR8",2011,24.7,"Méditerranée"
"Y15-24","FR81",2011,29.8,"Languedoc-Roussillon"
"Y15-24","FR82",2011,22.9,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2011,NA,"Corse"
"Y15-24","FRA",2011,56.2,"Départements d'outre-mer"
"Y15-24","FRA1",2011,53.2,"Guadeloupe"
"Y15-24","FRA2",2011,56.8,"Martinique"
"Y15-24","FRA3",2011,46.4,"Guyane"
"Y15-24","FRA4",2011,58.5,"La Réunion"
"Y15-24","HR",2011,36.7,"Croatia"
"Y15-24","HR0",2011,36.7,"Hrvatska"
"Y15-24","HR03",2011,32.9,"Jadranska Hrvatska"
"Y15-24","HR04",2011,38.3,"Kontinentalna Hrvatska"
"Y15-24","HU",2011,26,"Hungary"
"Y15-24","HU1",2011,20.2,"Közép-Magyarország"
"Y15-24","HU10",2011,20.2,"Közép-Magyarország"
"Y15-24","HU2",2011,22,"Dunántúl"
"Y15-24","HU21",2011,21.2,"Közép-Dunántúl"
"Y15-24","HU22",2011,17.4,"Nyugat-Dunántúl"
"Y15-24","HU23",2011,28.7,"Dél-Dunántúl"
"Y15-24","HU3",2011,32.3,"Alföld és Észak"
"Y15-24","HU31",2011,35.8,"Észak-Magyarország"
"Y15-24","HU32",2011,33.4,"Észak-Alföld"
"Y15-24","HU33",2011,27.3,"Dél-Alföld"
"Y15-24","IE",2011,29.1,"Ireland"
"Y15-24","IE0",2011,29.1,"Éire/Ireland"
"Y15-24","IE01",2011,32.8,"Border, Midland and Western"
"Y15-24","IE02",2011,27.8,"Southern and Eastern"
"Y15-24","IS",2011,14.4,"Iceland"
"Y15-24","IS0",2011,14.4,"Ísland"
"Y15-24","IS00",2011,14.4,"Ísland"
"Y15-24","IT",2011,29.2,"Italy"
"Y15-24","ITC",2011,22.4,"Nord-Ovest"
"Y15-24","ITC1",2011,25,"Piemonte"
"Y15-24","ITC2",2011,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2011,25.9,"Liguria"
"Y15-24","ITC4",2011,20.8,"Lombardia"
"Y15-24","ITF",2011,39.4,"Sud"
"Y15-24","ITF1",2011,26.5,"Abruzzo"
"Y15-24","ITF2",2011,29.3,"Molise"
"Y15-24","ITF3",2011,44.6,"Campania"
"Y15-24","ITF4",2011,37.5,"Puglia"
"Y15-24","ITF5",2011,39.7,"Basilicata"
"Y15-24","ITF6",2011,39.8,"Calabria"
"Y15-24","ITG",2011,42.4,"Isole"
"Y15-24","ITG1",2011,42.5,"Sicilia"
"Y15-24","ITG2",2011,42.2,"Sardegna"
"Y15-24","ITH",2011,19.5,"Nord-Est"
"Y15-24","ITH1",2011,9.1,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2011,14.4,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2011,19.7,"Veneto"
"Y15-24","ITH4",2011,21,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2011,21.8,"Emilia-Romagna"
"Y15-24","ITI",2011,28.6,"Centro (IT)"
"Y15-24","ITI1",2011,24.3,"Toscana"
"Y15-24","ITI2",2011,22.6,"Umbria"
"Y15-24","ITI3",2011,23.8,"Marche"
"Y15-24","ITI4",2011,33.8,"Lazio"
"Y15-24","LT",2011,32.6,"Lithuania"
"Y15-24","LT0",2011,32.6,"Lietuva"
"Y15-24","LT00",2011,32.6,"Lietuva"
"Y15-24","LU",2011,16.8,"Luxembourg"
"Y15-24","LU0",2011,16.8,"Luxembourg"
"Y15-24","LU00",2011,16.8,"Luxembourg"
"Y15-24","LV",2011,31,"Latvia"
"Y15-24","LV0",2011,31,"Latvija"
"Y15-24","LV00",2011,31,"Latvija"
"Y15-24","MK",2011,55.3,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2011,55.3,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2011,55.3,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2011,13.3,"Malta"
"Y15-24","MT0",2011,13.3,"Malta"
"Y15-24","MT00",2011,13.3,"Malta"
"Y15-24","NL",2011,10,"Netherlands"
"Y15-24","NL1",2011,11.8,"Noord-Nederland"
"Y15-24","NL11",2011,12.7,"Groningen"
"Y15-24","NL12",2011,10.8,"Friesland (NL)"
"Y15-24","NL13",2011,11.8,"Drenthe"
"Y15-24","NL2",2011,9.4,"Oost-Nederland"
"Y15-24","NL21",2011,10.3,"Overijssel"
"Y15-24","NL22",2011,8.9,"Gelderland"
"Y15-24","NL23",2011,9.3,"Flevoland"
"Y15-24","NL3",2011,10.2,"West-Nederland"
"Y15-24","NL31",2011,8.4,"Utrecht"
"Y15-24","NL32",2011,10.8,"Noord-Holland"
"Y15-24","NL33",2011,10.8,"Zuid-Holland"
"Y15-24","NL34",2011,5.4,"Zeeland"
"Y15-24","NL4",2011,9.4,"Zuid-Nederland"
"Y15-24","NL41",2011,9.2,"Noord-Brabant"
"Y15-24","NL42",2011,9.9,"Limburg (NL)"
"Y15-24","NO",2011,8.7,"Norway"
"Y15-24","NO0",2011,8.7,"Norge"
"Y15-24","NO01",2011,9.6,"Oslo og Akershus"
"Y15-24","NO02",2011,6.4,"Hedmark og Oppland"
"Y15-24","NO03",2011,9,"Sør-Østlandet"
"Y15-24","NO04",2011,6.6,"Agder og Rogaland"
"Y15-24","NO05",2011,8.4,"Vestlandet"
"Y15-24","NO06",2011,9.7,"Trøndelag"
"Y15-24","NO07",2011,10.2,"Nord-Norge"
"Y15-24","PL",2011,25.8,"Poland"
"Y15-24","PL1",2011,23,"Region Centralny"
"Y15-24","PL11",2011,23.6,"Lódzkie"
"Y15-24","PL12",2011,22.6,"Mazowieckie"
"Y15-24","PL2",2011,23.6,"Region Poludniowy"
"Y15-24","PL21",2011,22.9,"Malopolskie"
"Y15-24","PL22",2011,24.2,"Slaskie"
"Y15-24","PL3",2011,32.7,"Region Wschodni"
"Y15-24","PL31",2011,31.9,"Lubelskie"
"Y15-24","PL32",2011,36.6,"Podkarpackie"
"Y15-24","PL33",2011,34.4,"Swietokrzyskie"
"Y15-24","PL34",2011,25,"Podlaskie"
"Y15-24","PL4",2011,25.6,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2011,23.3,"Wielkopolskie"
"Y15-24","PL42",2011,32.9,"Zachodniopomorskie"
"Y15-24","PL43",2011,25.7,"Lubuskie"
"Y15-24","PL5",2011,23.7,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2011,24.5,"Dolnoslaskie"
"Y15-24","PL52",2011,21.3,"Opolskie"
"Y15-24","PL6",2011,25.6,"Region Pólnocny"
"Y15-24","PL61",2011,28.3,"Kujawsko-Pomorskie"
"Y15-24","PL62",2011,27.6,"Warminsko-Mazurskie"
"Y15-24","PL63",2011,22,"Pomorskie"
"Y15-24","PT",2011,30.3,"Portugal"
"Y15-24","PT1",2011,30,"Continente"
"Y15-24","PT11",2011,29,"Norte"
"Y15-24","PT15",2011,37,"Algarve"
"Y15-24","PT16",2011,26.4,"Centro (PT)"
"Y15-24","PT17",2011,32.6,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2011,32.7,"Alentejo"
"Y15-24","PT2",2011,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2011,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2011,39.4,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2011,39.4,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2011,23.9,"Romania"
"Y15-24","RO1",2011,27.6,"Macroregiunea unu"
"Y15-24","RO11",2011,20.9,"Nord-Vest"
"Y15-24","RO12",2011,35.8,"Centru"
"Y15-24","RO2",2011,19,"Macroregiunea doi"
"Y15-24","RO21",2011,12.2,"Nord-Est"
"Y15-24","RO22",2011,30.7,"Sud-Est"
"Y15-24","RO3",2011,28.7,"Macroregiunea trei"
"Y15-24","RO31",2011,32.9,"Sud - Muntenia"
"Y15-24","RO32",2011,22.1,"Bucuresti - Ilfov"
"Y15-24","RO4",2011,20.1,"Macroregiunea patru"
"Y15-24","RO41",2011,19.3,"Sud-Vest Oltenia"
"Y15-24","RO42",2011,21,"Vest"
"Y15-24","SE",2011,22.8,"Sweden"
"Y15-24","SE1",2011,21.5,"Östra Sverige"
"Y15-24","SE11",2011,19.9,"Stockholm"
"Y15-24","SE12",2011,23.4,"Östra Mellansverige"
"Y15-24","SE2",2011,22.8,"Södra Sverige"
"Y15-24","SE21",2011,20.4,"Småland med öarna"
"Y15-24","SE22",2011,25.1,"Sydsverige"
"Y15-24","SE23",2011,22.1,"Västsverige"
"Y15-24","SE3",2011,25.6,"Norra Sverige"
"Y15-24","SE31",2011,24.5,"Norra Mellansverige"
"Y15-24","SE32",2011,29.3,"Mellersta Norrland"
"Y15-24","SE33",2011,24.7,"Övre Norrland"
"Y15-24","SI",2011,15.7,"Slovenia"
"Y15-24","SI0",2011,15.7,"Slovenija"
"Y15-24","SI03",2011,18,"Vzhodna Slovenija"
"Y15-24","SI04",2011,13.2,"Zahodna Slovenija"
"Y15-24","SK",2011,33.4,"Slovakia"
"Y15-24","SK0",2011,33.4,"Slovensko"
"Y15-24","SK01",2011,17,"Bratislavský kraj"
"Y15-24","SK02",2011,26.8,"Západné Slovensko"
"Y15-24","SK03",2011,36,"Stredné Slovensko"
"Y15-24","SK04",2011,42.2,"Východné Slovensko"
"Y15-24","TR",2011,16.7,"Turkey"
"Y15-24","TR1",2011,18.2,"Istanbul"
"Y15-24","TR10",2011,18.2,"Istanbul"
"Y15-24","TR2",2011,14.9,"Bati Marmara"
"Y15-24","TR21",2011,17.6,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2011,11.4,"Balikesir, Çanakkale"
"Y15-24","TR3",2011,19.2,"Ege"
"Y15-24","TR31",2011,25.5,"Izmir"
"Y15-24","TR32",2011,16.3,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2011,11.5,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2011,16.1,"Dogu Marmara"
"Y15-24","TR41",2011,12.9,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2011,19.4,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2011,16.9,"Bati Anadolu"
"Y15-24","TR51",2011,20.7,"Ankara"
"Y15-24","TR52",2011,11.2,"Konya, Karaman"
"Y15-24","TR6",2011,16.8,"Akdeniz"
"Y15-24","TR61",2011,16.4,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2011,16.3,"Adana, Mersin"
"Y15-24","TR63",2011,17.9,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2011,17,"Orta Anadolu"
"Y15-24","TR71",2011,14.1,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2011,18.7,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2011,12,"Bati Karadeniz"
"Y15-24","TR81",2011,20.7,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2011,9.8,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2011,9.6,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2011,18.8,"Dogu Karadeniz"
"Y15-24","TR90",2011,18.8,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2011,13.1,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2011,11.8,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2011,14.2,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2011,15.7,"Ortadogu Anadolu"
"Y15-24","TRB1",2011,17.2,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2011,14.6,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2011,15.4,"Güneydogu Anadolu"
"Y15-24","TRC1",2011,20.7,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2011,9.5,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2011,16.2,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2011,21.3,"United Kingdom"
"Y15-24","UKC",2011,22.1,"North East (UK)"
"Y15-24","UKC1",2011,23.6,"Tees Valley and Durham"
"Y15-24","UKC2",2011,20.9,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2011,24.2,"North West (UK)"
"Y15-24","UKD1",2011,23.5,"Cumbria"
"Y15-24","UKD3",2011,25.8,"Greater Manchester"
"Y15-24","UKD4",2011,22.3,"Lancashire"
"Y15-24","UKD6",2011,17.2,"Cheshire"
"Y15-24","UKD7",2011,27.1,"Merseyside"
"Y15-24","UKE",2011,23.9,"Yorkshire and The Humber"
"Y15-24","UKE1",2011,22,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2011,21.7,"North Yorkshire"
"Y15-24","UKE3",2011,27.1,"South Yorkshire"
"Y15-24","UKE4",2011,23.1,"West Yorkshire"
"Y15-24","UKF",2011,21,"East Midlands (UK)"
"Y15-24","UKF1",2011,24,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2011,19.8,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2011,15.7,"Lincolnshire"
"Y15-24","UKG",2011,24.2,"West Midlands (UK)"
"Y15-24","UKG1",2011,20.2,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2011,20,"Shropshire and Staffordshire"
"Y15-24","UKG3",2011,28.2,"West Midlands"
"Y15-24","UKH",2011,17.8,"East of England"
"Y15-24","UKH1",2011,16.2,"East Anglia"
"Y15-24","UKH2",2011,18.2,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2011,19.8,"Essex"
"Y15-24","UKI",2011,24.7,"London"
"Y15-24","UKI3",2011,25.5,"Inner London - West"
"Y15-24","UKI4",2011,31.5,"Inner London - East"
"Y15-24","UKI5",2011,25.5,"Outer London - East and North East"
"Y15-24","UKI6",2011,21.1,"Outer London - South"
"Y15-24","UKI7",2011,18.1,"Outer London - West and North West"
"Y15-24","UKJ",2011,16.1,"South East (UK)"
"Y15-24","UKJ1",2011,12.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2011,14.9,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2011,15.2,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2011,22.2,"Kent"
"Y15-24","UKK",2011,16.6,"South West (UK)"
"Y15-24","UKK1",2011,18.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2011,12.7,"Dorset and Somerset"
"Y15-24","UKK3",2011,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2011,19,"Devon"
"Y15-24","UKL",2011,25.3,"Wales"
"Y15-24","UKL1",2011,28.5,"West Wales and The Valleys"
"Y15-24","UKL2",2011,20.6,"East Wales"
"Y15-24","UKM",2011,21.7,"Scotland"
"Y15-24","UKM2",2011,20.9,"Eastern Scotland"
"Y15-24","UKM3",2011,26.2,"South Western Scotland"
"Y15-24","UKM5",2011,12.3,"North Eastern Scotland"
"Y15-24","UKM6",2011,15.5,"Highlands and Islands"
"Y15-24","UKN",2011,19.8,"Northern Ireland (UK)"
"Y15-24","UKN0",2011,19.8,"Northern Ireland (UK)"
"Y20-64","AT",2011,4.3,"Austria"
"Y20-64","AT1",2011,5.7,"Ostösterreich"
"Y20-64","AT11",2011,3.5,"Burgenland (AT)"
"Y20-64","AT12",2011,4.3,"Niederösterreich"
"Y20-64","AT13",2011,7.5,"Wien"
"Y20-64","AT2",2011,3.7,"Südösterreich"
"Y20-64","AT21",2011,4,"Kärnten"
"Y20-64","AT22",2011,3.6,"Steiermark"
"Y20-64","AT3",2011,3,"Westösterreich"
"Y20-64","AT31",2011,3.2,"Oberösterreich"
"Y20-64","AT32",2011,2.7,"Salzburg"
"Y20-64","AT33",2011,2.5,"Tirol"
"Y20-64","AT34",2011,3.7,"Vorarlberg"
"Y20-64","BE",2011,6.9,"Belgium"
"Y20-64","BE1",2011,16.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2011,16.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2011,4,"Vlaams Gewest"
"Y20-64","BE21",2011,5.5,"Prov. Antwerpen"
"Y20-64","BE22",2011,4.2,"Prov. Limburg (BE)"
"Y20-64","BE23",2011,3.5,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2011,3.4,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2011,3,"Prov. West-Vlaanderen"
"Y20-64","BE3",2011,9.2,"Région wallonne"
"Y20-64","BE31",2011,6.4,"Prov. Brabant Wallon"
"Y20-64","BE32",2011,11.3,"Prov. Hainaut"
"Y20-64","BE33",2011,9.3,"Prov. Liège"
"Y20-64","BE34",2011,6,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2011,7.6,"Prov. Namur"
"Y20-64","BG",2011,11,"Bulgaria"
"Y20-64","BG3",2011,12.8,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2011,12.5,"Severozapaden"
"Y20-64","BG32",2011,12.5,"Severen tsentralen"
"Y20-64","BG33",2011,15.2,"Severoiztochen"
"Y20-64","BG34",2011,11.2,"Yugoiztochen"
"Y20-64","BG4",2011,9.3,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2011,7.3,"Yugozapaden"
"Y20-64","BG42",2011,12.7,"Yuzhen tsentralen"
"Y20-64","CH",2011,3.9,"Switzerland"
"Y20-64","CH0",2011,3.9,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2011,6,"Région lémanique"
"Y20-64","CH02",2011,3.3,"Espace Mittelland"
"Y20-64","CH03",2011,4,"Nordwestschweiz"
"Y20-64","CH04",2011,3.6,"Zürich"
"Y20-64","CH05",2011,3.1,"Ostschweiz"
"Y20-64","CH06",2011,2.3,"Zentralschweiz"
"Y20-64","CH07",2011,5.8,"Ticino"
"Y20-64","CY",2011,7.8,"Cyprus"
"Y20-64","CY0",2011,7.8,"Kypros"
"Y20-64","CY00",2011,7.8,"Kypros"
"Y20-64","CZ",2011,6.5,"Czech Republic"
"Y20-64","CZ0",2011,6.5,"Ceská republika"
"Y20-64","CZ01",2011,3.5,"Praha"
"Y20-64","CZ02",2011,4.9,"Strední Cechy"
"Y20-64","CZ03",2011,5.2,"Jihozápad"
"Y20-64","CZ04",2011,9.1,"Severozápad"
"Y20-64","CZ05",2011,6.4,"Severovýchod"
"Y20-64","CZ06",2011,7,"Jihovýchod"
"Y20-64","CZ07",2011,7.4,"Strední Morava"
"Y20-64","CZ08",2011,9.2,"Moravskoslezsko"
"Y20-64","DE",2011,5.8,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2011,3.5,"Baden-Württemberg"
"Y20-64","DE11",2011,3.6,"Stuttgart"
"Y20-64","DE12",2011,4.1,"Karlsruhe"
"Y20-64","DE13",2011,2.9,"Freiburg"
"Y20-64","DE14",2011,3.1,"Tübingen"
"Y20-64","DE2",2011,3.2,"Bayern"
"Y20-64","DE21",2011,2.7,"Oberbayern"
"Y20-64","DE22",2011,2.7,"Niederbayern"
"Y20-64","DE23",2011,3.3,"Oberpfalz"
"Y20-64","DE24",2011,4.2,"Oberfranken"
"Y20-64","DE25",2011,3.9,"Mittelfranken"
"Y20-64","DE26",2011,3.4,"Unterfranken"
"Y20-64","DE27",2011,3.3,"Schwaben"
"Y20-64","DE3",2011,11.7,"Berlin"
"Y20-64","DE30",2011,11.7,"Berlin"
"Y20-64","DE4",2011,8.8,"Brandenburg"
"Y20-64","DE40",2011,8.8,"Brandenburg"
"Y20-64","DE5",2011,7.7,"Bremen"
"Y20-64","DE50",2011,7.7,"Bremen"
"Y20-64","DE6",2011,5.4,"Hamburg"
"Y20-64","DE60",2011,5.4,"Hamburg"
"Y20-64","DE7",2011,4.6,"Hessen"
"Y20-64","DE71",2011,4.5,"Darmstadt"
"Y20-64","DE72",2011,5,"Gießen"
"Y20-64","DE73",2011,4.5,"Kassel"
"Y20-64","DE8",2011,10.1,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2011,10.1,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2011,5.4,"Niedersachsen"
"Y20-64","DE91",2011,6.1,"Braunschweig"
"Y20-64","DE92",2011,6.5,"Hannover"
"Y20-64","DE93",2011,5.2,"Lüneburg"
"Y20-64","DE94",2011,4.1,"Weser-Ems"
"Y20-64","DEA",2011,6.2,"Nordrhein-Westfalen"
"Y20-64","DEA1",2011,6.7,"Düsseldorf"
"Y20-64","DEA2",2011,5.8,"Köln"
"Y20-64","DEA3",2011,5.3,"Münster"
"Y20-64","DEA4",2011,5.4,"Detmold"
"Y20-64","DEA5",2011,7.1,"Arnsberg"
"Y20-64","DEB",2011,4.6,"Rheinland-Pfalz"
"Y20-64","DEB1",2011,4.3,"Koblenz"
"Y20-64","DEB2",2011,4,"Trier"
"Y20-64","DEB3",2011,4.9,"Rheinhessen-Pfalz"
"Y20-64","DEC",2011,5.6,"Saarland"
"Y20-64","DEC0",2011,5.6,"Saarland"
"Y20-64","DED",2011,9.4,"Sachsen"
"Y20-64","DED2",2011,8.8,"Dresden"
"Y20-64","DED4",2011,9,"Chemnitz"
"Y20-64","DED5",2011,11.1,"Leipzig"
"Y20-64","DEE",2011,10.5,"Sachsen-Anhalt"
"Y20-64","DEE0",2011,10.5,"Sachsen-Anhalt"
"Y20-64","DEF",2011,5.7,"Schleswig-Holstein"
"Y20-64","DEF0",2011,5.7,"Schleswig-Holstein"
"Y20-64","DEG",2011,7.5,"Thüringen"
"Y20-64","DEG0",2011,7.5,"Thüringen"
"Y20-64","DK",2011,7,"Denmark"
"Y20-64","DK0",2011,7,"Danmark"
"Y20-64","DK01",2011,7.5,"Hovedstaden"
"Y20-64","DK02",2011,6.5,"Sjælland"
"Y20-64","DK03",2011,7.1,"Syddanmark"
"Y20-64","DK04",2011,6.2,"Midtjylland"
"Y20-64","DK05",2011,7.5,"Nordjylland"
"Y20-64","EA17",2011,9.9,"Euro area (17 countries)"
"Y20-64","EA18",2011,9.9,"Euro area (18 countries)"
"Y20-64","EA19",2011,10,"Euro area (19 countries)"
"Y20-64","EE",2011,12.2,"Estonia"
"Y20-64","EE0",2011,12.2,"Eesti"
"Y20-64","EE00",2011,12.2,"Eesti"
"Y20-64","EL",2011,17.8,"Greece"
"Y20-64","EL3",2011,17.9,"Attiki"
"Y20-64","EL30",2011,17.9,"Attiki"
"Y20-64","EL4",2011,15.3,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2011,14.4,"Voreio Aigaio"
"Y20-64","EL42",2011,14.9,"Notio Aigaio"
"Y20-64","EL43",2011,15.8,"Kriti"
"Y20-64","EL5",2011,19.6,"Voreia Ellada"
"Y20-64","EL51",2011,19.7,"Anatoliki Makedonia, Thraki"
"Y20-64","EL52",2011,19.6,"Kentriki Makedonia"
"Y20-64","EL53",2011,23.2,"Dytiki Makedonia"
"Y20-64","EL54",2011,16.5,"Ipeiros"
"Y20-64","EL6",2011,16.6,"Kentriki Ellada"
"Y20-64","EL61",2011,16.8,"Thessalia"
"Y20-64","EL62",2011,14.2,"Ionia Nisia"
"Y20-64","EL63",2011,17.3,"Dytiki Ellada"
"Y20-64","EL64",2011,19,"Sterea Ellada"
"Y20-64","EL65",2011,13.9,"Peloponnisos"
"Y20-64","ES",2011,20.9,"Spain"
"Y20-64","ES1",2011,16.9,"Noroeste (ES)"
"Y20-64","ES11",2011,17,"Galicia"
"Y20-64","ES12",2011,17.6,"Principado de Asturias"
"Y20-64","ES13",2011,15.1,"Cantabria"
"Y20-64","ES2",2011,13.9,"Noreste (ES)"
"Y20-64","ES21",2011,12.2,"País Vasco"
"Y20-64","ES22",2011,12.6,"Comunidad Foral de Navarra"
"Y20-64","ES23",2011,16.4,"La Rioja"
"Y20-64","ES24",2011,16.6,"Aragón"
"Y20-64","ES3",2011,15.9,"Comunidad de Madrid"
"Y20-64","ES30",2011,15.9,"Comunidad de Madrid"
"Y20-64","ES4",2011,20.2,"Centro (ES)"
"Y20-64","ES41",2011,16.5,"Castilla y León"
"Y20-64","ES42",2011,22.5,"Castilla-la Mancha"
"Y20-64","ES43",2011,24.4,"Extremadura"
"Y20-64","ES5",2011,20.5,"Este (ES)"
"Y20-64","ES51",2011,18.6,"Cataluña"
"Y20-64","ES52",2011,23.4,"Comunidad Valenciana"
"Y20-64","ES53",2011,21.3,"Illes Balears"
"Y20-64","ES6",2011,28.6,"Sur (ES)"
"Y20-64","ES61",2011,29.5,"Andalucía"
"Y20-64","ES62",2011,24.2,"Región de Murcia"
"Y20-64","ES63",2011,26,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2011,21.5,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2011,28.9,"Canarias (ES)"
"Y20-64","ES70",2011,28.9,"Canarias (ES)"
"Y20-64","EU15",2011,9.3,"European Union (15 countries)"
"Y20-64","EU27",2011,9.3,"European Union (27 countries)"
"Y20-64","EU28",2011,9.4,"European Union (28 countries)"
"Y20-64","FI",2011,7.1,"Finland"
"Y20-64","FI1",2011,7.1,"Manner-Suomi"
"Y20-64","FI19",2011,7.5,"Länsi-Suomi"
"Y20-64","FI1B",2011,5.2,"Helsinki-Uusimaa"
"Y20-64","FI1C",2011,7.8,"Etelä-Suomi"
"Y20-64","FI1D",2011,8.7,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2011,NA,"Åland"
"Y20-64","FI20",2011,NA,"Åland"
"Y20-64","FR",2011,8.9,"France"
"Y20-64","FR1",2011,8,"Île de France"
"Y20-64","FR10",2011,8,"Île de France"
"Y20-64","FR2",2011,8.5,"Bassin Parisien"
"Y20-64","FR21",2011,9.7,"Champagne-Ardenne"
"Y20-64","FR22",2011,8.5,"Picardie"
"Y20-64","FR23",2011,8.5,"Haute-Normandie"
"Y20-64","FR24",2011,8,"Centre (FR)"
"Y20-64","FR25",2011,8.9,"Basse-Normandie"
"Y20-64","FR26",2011,8.3,"Bourgogne"
"Y20-64","FR3",2011,11.5,"Nord - Pas-de-Calais"
"Y20-64","FR30",2011,11.5,"Nord - Pas-de-Calais"
"Y20-64","FR4",2011,8.3,"Est (FR)"
"Y20-64","FR41",2011,9.9,"Lorraine"
"Y20-64","FR42",2011,6.8,"Alsace"
"Y20-64","FR43",2011,7.6,"Franche-Comté"
"Y20-64","FR5",2011,7.5,"Ouest (FR)"
"Y20-64","FR51",2011,8.1,"Pays de la Loire"
"Y20-64","FR52",2011,6.8,"Bretagne"
"Y20-64","FR53",2011,7.6,"Poitou-Charentes"
"Y20-64","FR6",2011,8.2,"Sud-Ouest (FR)"
"Y20-64","FR61",2011,8.6,"Aquitaine"
"Y20-64","FR62",2011,7.9,"Midi-Pyrénées"
"Y20-64","FR63",2011,7.4,"Limousin"
"Y20-64","FR7",2011,7.5,"Centre-Est (FR)"
"Y20-64","FR71",2011,7.4,"Rhône-Alpes"
"Y20-64","FR72",2011,8,"Auvergne"
"Y20-64","FR8",2011,9.9,"Méditerranée"
"Y20-64","FR81",2011,11.3,"Languedoc-Roussillon"
"Y20-64","FR82",2011,9.4,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2011,NA,"Corse"
"Y20-64","FRA",2011,24.7,"Départements d'outre-mer"
"Y20-64","FRA1",2011,22.4,"Guadeloupe"
"Y20-64","FRA2",2011,20.6,"Martinique"
"Y20-64","FRA3",2011,20.6,"Guyane"
"Y20-64","FRA4",2011,28.7,"La Réunion"
"Y20-64","HR",2011,13.2,"Croatia"
"Y20-64","HR0",2011,13.2,"Hrvatska"
"Y20-64","HR03",2011,12.6,"Jadranska Hrvatska"
"Y20-64","HR04",2011,13.5,"Kontinentalna Hrvatska"
"Y20-64","HU",2011,11,"Hungary"
"Y20-64","HU1",2011,9,"Közép-Magyarország"
"Y20-64","HU10",2011,9,"Közép-Magyarország"
"Y20-64","HU2",2011,9.7,"Dunántúl"
"Y20-64","HU21",2011,9.3,"Közép-Dunántúl"
"Y20-64","HU22",2011,7.3,"Nyugat-Dunántúl"
"Y20-64","HU23",2011,12.9,"Dél-Dunántúl"
"Y20-64","HU3",2011,13.7,"Alföld és Észak"
"Y20-64","HU31",2011,16.3,"Észak-Magyarország"
"Y20-64","HU32",2011,14.5,"Észak-Alföld"
"Y20-64","HU33",2011,10.4,"Dél-Alföld"
"Y20-64","IE",2011,14.4,"Ireland"
"Y20-64","IE0",2011,14.4,"Éire/Ireland"
"Y20-64","IE01",2011,15.6,"Border, Midland and Western"
"Y20-64","IE02",2011,14,"Southern and Eastern"
"Y20-64","IS",2011,6.4,"Iceland"
"Y20-64","IS0",2011,6.4,"Ísland"
"Y20-64","IS00",2011,6.4,"Ísland"
"Y20-64","IT",2011,8.1,"Italy"
"Y20-64","ITC",2011,6,"Nord-Ovest"
"Y20-64","ITC1",2011,7.3,"Piemonte"
"Y20-64","ITC2",2011,5,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2011,6.1,"Liguria"
"Y20-64","ITC4",2011,5.4,"Lombardia"
"Y20-64","ITF",2011,13,"Sud"
"Y20-64","ITF1",2011,8.4,"Abruzzo"
"Y20-64","ITF2",2011,9.9,"Molise"
"Y20-64","ITF3",2011,15,"Campania"
"Y20-64","ITF4",2011,12.8,"Puglia"
"Y20-64","ITF5",2011,11.6,"Basilicata"
"Y20-64","ITF6",2011,12.4,"Calabria"
"Y20-64","ITG",2011,13.6,"Isole"
"Y20-64","ITG1",2011,13.8,"Sicilia"
"Y20-64","ITG2",2011,13.3,"Sardegna"
"Y20-64","ITH",2011,4.7,"Nord-Est"
"Y20-64","ITH1",2011,3,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2011,4.2,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2011,4.7,"Veneto"
"Y20-64","ITH4",2011,4.9,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2011,5,"Emilia-Romagna"
"Y20-64","ITI",2011,7.4,"Centro (IT)"
"Y20-64","ITI1",2011,6.2,"Toscana"
"Y20-64","ITI2",2011,6.2,"Umbria"
"Y20-64","ITI3",2011,6.7,"Marche"
"Y20-64","ITI4",2011,8.5,"Lazio"
"Y20-64","LT",2011,15.4,"Lithuania"
"Y20-64","LT0",2011,15.4,"Lietuva"
"Y20-64","LT00",2011,15.4,"Lietuva"
"Y20-64","LU",2011,4.8,"Luxembourg"
"Y20-64","LU0",2011,4.8,"Luxembourg"
"Y20-64","LU00",2011,4.8,"Luxembourg"
"Y20-64","LV",2011,16.1,"Latvia"
"Y20-64","LV0",2011,16.1,"Latvija"
"Y20-64","LV00",2011,16.1,"Latvija"
"Y20-64","MK",2011,31,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2011,31,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2011,31,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2011,5.6,"Malta"
"Y20-64","MT0",2011,5.6,"Malta"
"Y20-64","MT00",2011,5.6,"Malta"
"Y20-64","NL",2011,4.4,"Netherlands"
"Y20-64","NL1",2011,5.1,"Noord-Nederland"
"Y20-64","NL11",2011,6.3,"Groningen"
"Y20-64","NL12",2011,4.5,"Friesland (NL)"
"Y20-64","NL13",2011,4.6,"Drenthe"
"Y20-64","NL2",2011,4.1,"Oost-Nederland"
"Y20-64","NL21",2011,4.2,"Overijssel"
"Y20-64","NL22",2011,4,"Gelderland"
"Y20-64","NL23",2011,4.7,"Flevoland"
"Y20-64","NL3",2011,4.5,"West-Nederland"
"Y20-64","NL31",2011,3.9,"Utrecht"
"Y20-64","NL32",2011,4.4,"Noord-Holland"
"Y20-64","NL33",2011,5.1,"Zuid-Holland"
"Y20-64","NL34",2011,3,"Zeeland"
"Y20-64","NL4",2011,4.1,"Zuid-Nederland"
"Y20-64","NL41",2011,4.1,"Noord-Brabant"
"Y20-64","NL42",2011,4.2,"Limburg (NL)"
"Y20-64","NO",2011,2.9,"Norway"
"Y20-64","NO0",2011,2.9,"Norge"
"Y20-64","NO01",2011,3,"Oslo og Akershus"
"Y20-64","NO02",2011,2.7,"Hedmark og Oppland"
"Y20-64","NO03",2011,3.4,"Sør-Østlandet"
"Y20-64","NO04",2011,1.9,"Agder og Rogaland"
"Y20-64","NO05",2011,2.8,"Vestlandet"
"Y20-64","NO06",2011,3,"Trøndelag"
"Y20-64","NO07",2011,3,"Nord-Norge"
"Y20-64","PL",2011,9.5,"Poland"
"Y20-64","PL1",2011,8.2,"Region Centralny"
"Y20-64","PL11",2011,9.2,"Lódzkie"
"Y20-64","PL12",2011,7.7,"Mazowieckie"
"Y20-64","PL2",2011,9.2,"Region Poludniowy"
"Y20-64","PL21",2011,9.3,"Malopolskie"
"Y20-64","PL22",2011,9,"Slaskie"
"Y20-64","PL3",2011,11.3,"Region Wschodni"
"Y20-64","PL31",2011,10.3,"Lubelskie"
"Y20-64","PL32",2011,12.4,"Podkarpackie"
"Y20-64","PL33",2011,13.1,"Swietokrzyskie"
"Y20-64","PL34",2011,9.3,"Podlaskie"
"Y20-64","PL4",2011,9.4,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2011,8.5,"Wielkopolskie"
"Y20-64","PL42",2011,11.5,"Zachodniopomorskie"
"Y20-64","PL43",2011,9.3,"Lubuskie"
"Y20-64","PL5",2011,10.2,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2011,10.5,"Dolnoslaskie"
"Y20-64","PL52",2011,9.2,"Opolskie"
"Y20-64","PL6",2011,9.5,"Region Pólnocny"
"Y20-64","PL61",2011,10.8,"Kujawsko-Pomorskie"
"Y20-64","PL62",2011,9.3,"Warminsko-Mazurskie"
"Y20-64","PL63",2011,8.3,"Pomorskie"
"Y20-64","PT",2011,12.8,"Portugal"
"Y20-64","PT1",2011,12.8,"Continente"
"Y20-64","PT11",2011,13,"Norte"
"Y20-64","PT15",2011,15.6,"Algarve"
"Y20-64","PT16",2011,10.6,"Centro (PT)"
"Y20-64","PT17",2011,13.9,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2011,12.6,"Alentejo"
"Y20-64","PT2",2011,10.8,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2011,10.8,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2011,13.3,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2011,13.3,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2011,7.2,"Romania"
"Y20-64","RO1",2011,7.5,"Macroregiunea unu"
"Y20-64","RO11",2011,5,"Nord-Vest"
"Y20-64","RO12",2011,10.4,"Centru"
"Y20-64","RO2",2011,6.9,"Macroregiunea doi"
"Y20-64","RO21",2011,4.9,"Nord-Est"
"Y20-64","RO22",2011,9.6,"Sud-Est"
"Y20-64","RO3",2011,7.8,"Macroregiunea trei"
"Y20-64","RO31",2011,10,"Sud - Muntenia"
"Y20-64","RO32",2011,5.2,"Bucuresti - Ilfov"
"Y20-64","RO4",2011,6.3,"Macroregiunea patru"
"Y20-64","RO41",2011,7,"Sud-Vest Oltenia"
"Y20-64","RO42",2011,5.5,"Vest"
"Y20-64","SE",2011,6.9,"Sweden"
"Y20-64","SE1",2011,6.3,"Östra Sverige"
"Y20-64","SE11",2011,5.6,"Stockholm"
"Y20-64","SE12",2011,7.5,"Östra Mellansverige"
"Y20-64","SE2",2011,7.1,"Södra Sverige"
"Y20-64","SE21",2011,6.4,"Småland med öarna"
"Y20-64","SE22",2011,8.5,"Sydsverige"
"Y20-64","SE23",2011,6.5,"Västsverige"
"Y20-64","SE3",2011,7.4,"Norra Sverige"
"Y20-64","SE31",2011,7.6,"Norra Mellansverige"
"Y20-64","SE32",2011,7.6,"Mellersta Norrland"
"Y20-64","SE33",2011,7,"Övre Norrland"
"Y20-64","SI",2011,8.2,"Slovenia"
"Y20-64","SI0",2011,8.2,"Slovenija"
"Y20-64","SI03",2011,9.3,"Vzhodna Slovenija"
"Y20-64","SI04",2011,7,"Zahodna Slovenija"
"Y20-64","SK",2011,13.2,"Slovakia"
"Y20-64","SK0",2011,13.2,"Slovensko"
"Y20-64","SK01",2011,5.7,"Bratislavský kraj"
"Y20-64","SK02",2011,10.5,"Západné Slovensko"
"Y20-64","SK03",2011,15.2,"Stredné Slovensko"
"Y20-64","SK04",2011,18.1,"Východné Slovensko"
"Y20-64","TR",2011,8.6,"Turkey"
"Y20-64","TR1",2011,10.7,"Istanbul"
"Y20-64","TR10",2011,10.7,"Istanbul"
"Y20-64","TR2",2011,6.2,"Bati Marmara"
"Y20-64","TR21",2011,7.9,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2011,4.3,"Balikesir, Çanakkale"
"Y20-64","TR3",2011,9,"Ege"
"Y20-64","TR31",2011,13.3,"Izmir"
"Y20-64","TR32",2011,7.5,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2011,4.4,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2011,8.5,"Dogu Marmara"
"Y20-64","TR41",2011,6.5,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2011,10.5,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2011,7.4,"Bati Anadolu"
"Y20-64","TR51",2011,8.2,"Ankara"
"Y20-64","TR52",2011,5.6,"Konya, Karaman"
"Y20-64","TR6",2011,9.4,"Akdeniz"
"Y20-64","TR61",2011,8.5,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2011,9.3,"Adana, Mersin"
"Y20-64","TR63",2011,10.5,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2011,8.6,"Orta Anadolu"
"Y20-64","TR71",2011,7,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2011,9.7,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2011,5.5,"Bati Karadeniz"
"Y20-64","TR81",2011,7,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2011,5.7,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2011,4.8,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2011,5.5,"Dogu Karadeniz"
"Y20-64","TR90",2011,5.5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2011,7.3,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2011,5.7,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2011,8.8,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2011,9.2,"Ortadogu Anadolu"
"Y20-64","TRB1",2011,7.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2011,10.8,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2011,9.8,"Güneydogu Anadolu"
"Y20-64","TRC1",2011,12.7,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2011,6.8,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2011,9.8,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2011,7,"United Kingdom"
"Y20-64","UKC",2011,9.3,"North East (UK)"
"Y20-64","UKC1",2011,10.5,"Tees Valley and Durham"
"Y20-64","UKC2",2011,8.3,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2011,7.2,"North West (UK)"
"Y20-64","UKD1",2011,6.1,"Cumbria"
"Y20-64","UKD3",2011,8.4,"Greater Manchester"
"Y20-64","UKD4",2011,5.6,"Lancashire"
"Y20-64","UKD6",2011,4.7,"Cheshire"
"Y20-64","UKD7",2011,8.6,"Merseyside"
"Y20-64","UKE",2011,8.2,"Yorkshire and The Humber"
"Y20-64","UKE1",2011,8.4,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2011,6,"North Yorkshire"
"Y20-64","UKE3",2011,9.1,"South Yorkshire"
"Y20-64","UKE4",2011,8.5,"West Yorkshire"
"Y20-64","UKF",2011,6.5,"East Midlands (UK)"
"Y20-64","UKF1",2011,7.1,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2011,6.2,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2011,5.8,"Lincolnshire"
"Y20-64","UKG",2011,7.9,"West Midlands (UK)"
"Y20-64","UKG1",2011,5.1,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2011,6.8,"Shropshire and Staffordshire"
"Y20-64","UKG3",2011,10.1,"West Midlands"
"Y20-64","UKH",2011,5.8,"East of England"
"Y20-64","UKH1",2011,5.7,"East Anglia"
"Y20-64","UKH2",2011,5.8,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2011,6.1,"Essex"
"Y20-64","UKI",2011,9,"London"
"Y20-64","UKI3",2011,7,"Inner London - West"
"Y20-64","UKI4",2011,11,"Inner London - East"
"Y20-64","UKI5",2011,10.1,"Outer London - East and North East"
"Y20-64","UKI6",2011,7.3,"Outer London - South"
"Y20-64","UKI7",2011,7.7,"Outer London - West and North West"
"Y20-64","UKJ",2011,5.2,"South East (UK)"
"Y20-64","UKJ1",2011,4.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2011,4.6,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2011,5.2,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2011,7.1,"Kent"
"Y20-64","UKK",2011,5.7,"South West (UK)"
"Y20-64","UKK1",2011,5.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2011,5.6,"Dorset and Somerset"
"Y20-64","UKK3",2011,5.8,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2011,5.6,"Devon"
"Y20-64","UKL",2011,7.3,"Wales"
"Y20-64","UKL1",2011,8.6,"West Wales and The Valleys"
"Y20-64","UKL2",2011,5,"East Wales"
"Y20-64","UKM",2011,6.8,"Scotland"
"Y20-64","UKM2",2011,6.1,"Eastern Scotland"
"Y20-64","UKM3",2011,8.4,"South Western Scotland"
"Y20-64","UKM5",2011,4,"North Eastern Scotland"
"Y20-64","UKM6",2011,6.3,"Highlands and Islands"
"Y20-64","UKN",2011,6.5,"Northern Ireland (UK)"
"Y20-64","UKN0",2011,6.5,"Northern Ireland (UK)"
"Y_GE15","AT",2011,4.6,"Austria"
"Y_GE15","AT1",2011,6.1,"Ostösterreich"
"Y_GE15","AT11",2011,3.8,"Burgenland (AT)"
"Y_GE15","AT12",2011,4.5,"Niederösterreich"
"Y_GE15","AT13",2011,8,"Wien"
"Y_GE15","AT2",2011,3.8,"Südösterreich"
"Y_GE15","AT21",2011,4.3,"Kärnten"
"Y_GE15","AT22",2011,3.6,"Steiermark"
"Y_GE15","AT3",2011,3.2,"Westösterreich"
"Y_GE15","AT31",2011,3.4,"Oberösterreich"
"Y_GE15","AT32",2011,2.9,"Salzburg"
"Y_GE15","AT33",2011,2.7,"Tirol"
"Y_GE15","AT34",2011,4.1,"Vorarlberg"
"Y_GE15","BE",2011,7.1,"Belgium"
"Y_GE15","BE1",2011,16.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2011,16.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2011,4.3,"Vlaams Gewest"
"Y_GE15","BE21",2011,5.7,"Prov. Antwerpen"
"Y_GE15","BE22",2011,4.6,"Prov. Limburg (BE)"
"Y_GE15","BE23",2011,3.8,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2011,3.5,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2011,3.2,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2011,9.5,"Région wallonne"
"Y_GE15","BE31",2011,6.7,"Prov. Brabant Wallon"
"Y_GE15","BE32",2011,11.7,"Prov. Hainaut"
"Y_GE15","BE33",2011,9.5,"Prov. Liège"
"Y_GE15","BE34",2011,6.2,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2011,8,"Prov. Namur"
"Y_GE15","BG",2011,11.3,"Bulgaria"
"Y_GE15","BG3",2011,13.1,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2011,12.8,"Severozapaden"
"Y_GE15","BG32",2011,12.8,"Severen tsentralen"
"Y_GE15","BG33",2011,15.4,"Severoiztochen"
"Y_GE15","BG34",2011,11.5,"Yugoiztochen"
"Y_GE15","BG4",2011,9.5,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2011,7.5,"Yugozapaden"
"Y_GE15","BG42",2011,12.9,"Yuzhen tsentralen"
"Y_GE15","CH",2011,4,"Switzerland"
"Y_GE15","CH0",2011,4,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2011,6.2,"Région lémanique"
"Y_GE15","CH02",2011,3.5,"Espace Mittelland"
"Y_GE15","CH03",2011,4.1,"Nordwestschweiz"
"Y_GE15","CH04",2011,3.6,"Zürich"
"Y_GE15","CH05",2011,3.2,"Ostschweiz"
"Y_GE15","CH06",2011,2.4,"Zentralschweiz"
"Y_GE15","CH07",2011,6,"Ticino"
"Y_GE15","CY",2011,7.9,"Cyprus"
"Y_GE15","CY0",2011,7.9,"Kypros"
"Y_GE15","CY00",2011,7.9,"Kypros"
"Y_GE15","CZ",2011,6.7,"Czech Republic"
"Y_GE15","CZ0",2011,6.7,"Ceská republika"
"Y_GE15","CZ01",2011,3.6,"Praha"
"Y_GE15","CZ02",2011,5.1,"Strední Cechy"
"Y_GE15","CZ03",2011,5.3,"Jihozápad"
"Y_GE15","CZ04",2011,9.5,"Severozápad"
"Y_GE15","CZ05",2011,6.6,"Severovýchod"
"Y_GE15","CZ06",2011,7.2,"Jihovýchod"
"Y_GE15","CZ07",2011,7.6,"Strední Morava"
"Y_GE15","CZ08",2011,9.3,"Moravskoslezsko"
"Y_GE15","DE",2011,5.8,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2011,3.6,"Baden-Württemberg"
"Y_GE15","DE11",2011,3.6,"Stuttgart"
"Y_GE15","DE12",2011,4.2,"Karlsruhe"
"Y_GE15","DE13",2011,3,"Freiburg"
"Y_GE15","DE14",2011,3.1,"Tübingen"
"Y_GE15","DE2",2011,3.3,"Bayern"
"Y_GE15","DE21",2011,2.7,"Oberbayern"
"Y_GE15","DE22",2011,2.8,"Niederbayern"
"Y_GE15","DE23",2011,3.4,"Oberpfalz"
"Y_GE15","DE24",2011,4.2,"Oberfranken"
"Y_GE15","DE25",2011,4,"Mittelfranken"
"Y_GE15","DE26",2011,3.5,"Unterfranken"
"Y_GE15","DE27",2011,3.4,"Schwaben"
"Y_GE15","DE3",2011,11.6,"Berlin"
"Y_GE15","DE30",2011,11.6,"Berlin"
"Y_GE15","DE4",2011,8.8,"Brandenburg"
"Y_GE15","DE40",2011,8.8,"Brandenburg"
"Y_GE15","DE5",2011,7.7,"Bremen"
"Y_GE15","DE50",2011,7.7,"Bremen"
"Y_GE15","DE6",2011,5.3,"Hamburg"
"Y_GE15","DE60",2011,5.3,"Hamburg"
"Y_GE15","DE7",2011,4.7,"Hessen"
"Y_GE15","DE71",2011,4.7,"Darmstadt"
"Y_GE15","DE72",2011,5.1,"Gießen"
"Y_GE15","DE73",2011,4.4,"Kassel"
"Y_GE15","DE8",2011,10.1,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2011,10.1,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2011,5.5,"Niedersachsen"
"Y_GE15","DE91",2011,6.2,"Braunschweig"
"Y_GE15","DE92",2011,6.7,"Hannover"
"Y_GE15","DE93",2011,5.3,"Lüneburg"
"Y_GE15","DE94",2011,4.2,"Weser-Ems"
"Y_GE15","DEA",2011,6.3,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2011,6.7,"Düsseldorf"
"Y_GE15","DEA2",2011,6,"Köln"
"Y_GE15","DEA3",2011,5.3,"Münster"
"Y_GE15","DEA4",2011,5.5,"Detmold"
"Y_GE15","DEA5",2011,7.1,"Arnsberg"
"Y_GE15","DEB",2011,4.8,"Rheinland-Pfalz"
"Y_GE15","DEB1",2011,4.4,"Koblenz"
"Y_GE15","DEB2",2011,4.1,"Trier"
"Y_GE15","DEB3",2011,5.2,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2011,5.8,"Saarland"
"Y_GE15","DEC0",2011,5.8,"Saarland"
"Y_GE15","DED",2011,9.3,"Sachsen"
"Y_GE15","DED2",2011,8.6,"Dresden"
"Y_GE15","DED4",2011,8.8,"Chemnitz"
"Y_GE15","DED5",2011,11.1,"Leipzig"
"Y_GE15","DEE",2011,10.4,"Sachsen-Anhalt"
"Y_GE15","DEE0",2011,10.4,"Sachsen-Anhalt"
"Y_GE15","DEF",2011,5.8,"Schleswig-Holstein"
"Y_GE15","DEF0",2011,5.8,"Schleswig-Holstein"
"Y_GE15","DEG",2011,7.6,"Thüringen"
"Y_GE15","DEG0",2011,7.6,"Thüringen"
"Y_GE15","DK",2011,7.6,"Denmark"
"Y_GE15","DK0",2011,7.6,"Danmark"
"Y_GE15","DK01",2011,8.1,"Hovedstaden"
"Y_GE15","DK02",2011,7.2,"Sjælland"
"Y_GE15","DK03",2011,7.7,"Syddanmark"
"Y_GE15","DK04",2011,6.7,"Midtjylland"
"Y_GE15","DK05",2011,8,"Nordjylland"
"Y_GE15","EA17",2011,10.1,"Euro area (17 countries)"
"Y_GE15","EA18",2011,10.1,"Euro area (18 countries)"
"Y_GE15","EA19",2011,10.2,"Euro area (19 countries)"
"Y_GE15","EE",2011,12.3,"Estonia"
"Y_GE15","EE0",2011,12.3,"Eesti"
"Y_GE15","EE00",2011,12.3,"Eesti"
"Y_GE15","EL",2011,17.9,"Greece"
"Y_GE15","EL3",2011,18,"Attiki"
"Y_GE15","EL30",2011,18,"Attiki"
"Y_GE15","EL4",2011,15.5,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2011,15,"Voreio Aigaio"
"Y_GE15","EL42",2011,15.2,"Notio Aigaio"
"Y_GE15","EL43",2011,15.8,"Kriti"
"Y_GE15","EL5",2011,19.8,"Voreia Ellada"
"Y_GE15","EL51",2011,20.2,"Anatoliki Makedonia, Thraki"
"Y_GE15","EL52",2011,19.7,"Kentriki Makedonia"
"Y_GE15","EL53",2011,23.1,"Dytiki Makedonia"
"Y_GE15","EL54",2011,16.5,"Ipeiros"
"Y_GE15","EL6",2011,16.6,"Kentriki Ellada"
"Y_GE15","EL61",2011,16.8,"Thessalia"
"Y_GE15","EL62",2011,14.1,"Ionia Nisia"
"Y_GE15","EL63",2011,17.6,"Dytiki Ellada"
"Y_GE15","EL64",2011,19,"Sterea Ellada"
"Y_GE15","EL65",2011,13.8,"Peloponnisos"
"Y_GE15","ES",2011,21.4,"Spain"
"Y_GE15","ES1",2011,17.1,"Noroeste (ES)"
"Y_GE15","ES11",2011,17.3,"Galicia"
"Y_GE15","ES12",2011,17.8,"Principado de Asturias"
"Y_GE15","ES13",2011,15.3,"Cantabria"
"Y_GE15","ES2",2011,14.2,"Noreste (ES)"
"Y_GE15","ES21",2011,12.4,"País Vasco"
"Y_GE15","ES22",2011,13,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2011,17.2,"La Rioja"
"Y_GE15","ES24",2011,17.1,"Aragón"
"Y_GE15","ES3",2011,16.3,"Comunidad de Madrid"
"Y_GE15","ES30",2011,16.3,"Comunidad de Madrid"
"Y_GE15","ES4",2011,20.7,"Centro (ES)"
"Y_GE15","ES41",2011,16.9,"Castilla y León"
"Y_GE15","ES42",2011,23.1,"Castilla-la Mancha"
"Y_GE15","ES43",2011,25.1,"Extremadura"
"Y_GE15","ES5",2011,21.1,"Este (ES)"
"Y_GE15","ES51",2011,19.2,"Cataluña"
"Y_GE15","ES52",2011,24,"Comunidad Valenciana"
"Y_GE15","ES53",2011,21.9,"Illes Balears"
"Y_GE15","ES6",2011,29.3,"Sur (ES)"
"Y_GE15","ES61",2011,30.1,"Andalucía"
"Y_GE15","ES62",2011,25,"Región de Murcia"
"Y_GE15","ES63",2011,27.7,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2011,22.4,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2011,29.3,"Canarias (ES)"
"Y_GE15","ES70",2011,29.3,"Canarias (ES)"
"Y_GE15","EU15",2011,9.6,"European Union (15 countries)"
"Y_GE15","EU27",2011,9.6,"European Union (27 countries)"
"Y_GE15","EU28",2011,9.6,"European Union (28 countries)"
"Y_GE15","FI",2011,7.8,"Finland"
"Y_GE15","FI1",2011,7.8,"Manner-Suomi"
"Y_GE15","FI19",2011,8.3,"Länsi-Suomi"
"Y_GE15","FI1B",2011,5.8,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2011,8.5,"Etelä-Suomi"
"Y_GE15","FI1D",2011,9.4,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2011,NA,"Åland"
"Y_GE15","FI20",2011,NA,"Åland"
"Y_GE15","FR",2011,9.2,"France"
"Y_GE15","FR1",2011,8.2,"Île de France"
"Y_GE15","FR10",2011,8.2,"Île de France"
"Y_GE15","FR2",2011,9,"Bassin Parisien"
"Y_GE15","FR21",2011,10.3,"Champagne-Ardenne"
"Y_GE15","FR22",2011,9,"Picardie"
"Y_GE15","FR23",2011,8.9,"Haute-Normandie"
"Y_GE15","FR24",2011,8.3,"Centre (FR)"
"Y_GE15","FR25",2011,9.2,"Basse-Normandie"
"Y_GE15","FR26",2011,8.8,"Bourgogne"
"Y_GE15","FR3",2011,12.3,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2011,12.3,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2011,8.7,"Est (FR)"
"Y_GE15","FR41",2011,10.1,"Lorraine"
"Y_GE15","FR42",2011,7.4,"Alsace"
"Y_GE15","FR43",2011,7.9,"Franche-Comté"
"Y_GE15","FR5",2011,7.9,"Ouest (FR)"
"Y_GE15","FR51",2011,8.5,"Pays de la Loire"
"Y_GE15","FR52",2011,7.1,"Bretagne"
"Y_GE15","FR53",2011,8.1,"Poitou-Charentes"
"Y_GE15","FR6",2011,8.4,"Sud-Ouest (FR)"
"Y_GE15","FR61",2011,9,"Aquitaine"
"Y_GE15","FR62",2011,8.1,"Midi-Pyrénées"
"Y_GE15","FR63",2011,7.5,"Limousin"
"Y_GE15","FR7",2011,7.9,"Centre-Est (FR)"
"Y_GE15","FR71",2011,7.7,"Rhône-Alpes"
"Y_GE15","FR72",2011,8.4,"Auvergne"
"Y_GE15","FR8",2011,10.3,"Méditerranée"
"Y_GE15","FR81",2011,11.9,"Languedoc-Roussillon"
"Y_GE15","FR82",2011,9.7,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2011,NA,"Corse"
"Y_GE15","FRA",2011,25.3,"Départements d'outre-mer"
"Y_GE15","FRA1",2011,22.6,"Guadeloupe"
"Y_GE15","FRA2",2011,20.8,"Martinique"
"Y_GE15","FRA3",2011,21,"Guyane"
"Y_GE15","FRA4",2011,29.6,"La Réunion"
"Y_GE15","HR",2011,13.7,"Croatia"
"Y_GE15","HR0",2011,13.7,"Hrvatska"
"Y_GE15","HR03",2011,13.3,"Jadranska Hrvatska"
"Y_GE15","HR04",2011,13.9,"Kontinentalna Hrvatska"
"Y_GE15","HU",2011,11,"Hungary"
"Y_GE15","HU1",2011,9,"Közép-Magyarország"
"Y_GE15","HU10",2011,9,"Közép-Magyarország"
"Y_GE15","HU2",2011,9.7,"Dunántúl"
"Y_GE15","HU21",2011,9.5,"Közép-Dunántúl"
"Y_GE15","HU22",2011,7.3,"Nyugat-Dunántúl"
"Y_GE15","HU23",2011,12.9,"Dél-Dunántúl"
"Y_GE15","HU3",2011,13.8,"Alföld és Észak"
"Y_GE15","HU31",2011,16.4,"Észak-Magyarország"
"Y_GE15","HU32",2011,14.6,"Észak-Alföld"
"Y_GE15","HU33",2011,10.5,"Dél-Alföld"
"Y_GE15","IE",2011,14.6,"Ireland"
"Y_GE15","IE0",2011,14.6,"Éire/Ireland"
"Y_GE15","IE01",2011,15.9,"Border, Midland and Western"
"Y_GE15","IE02",2011,14.2,"Southern and Eastern"
"Y_GE15","IS",2011,7,"Iceland"
"Y_GE15","IS0",2011,7,"Ísland"
"Y_GE15","IS00",2011,7,"Ísland"
"Y_GE15","IT",2011,8.4,"Italy"
"Y_GE15","ITC",2011,6.3,"Nord-Ovest"
"Y_GE15","ITC1",2011,7.6,"Piemonte"
"Y_GE15","ITC2",2011,5.3,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2011,6.4,"Liguria"
"Y_GE15","ITC4",2011,5.7,"Lombardia"
"Y_GE15","ITF",2011,13.3,"Sud"
"Y_GE15","ITF1",2011,8.6,"Abruzzo"
"Y_GE15","ITF2",2011,9.9,"Molise"
"Y_GE15","ITF3",2011,15.4,"Campania"
"Y_GE15","ITF4",2011,13.2,"Puglia"
"Y_GE15","ITF5",2011,11.9,"Basilicata"
"Y_GE15","ITF6",2011,12.7,"Calabria"
"Y_GE15","ITG",2011,14,"Isole"
"Y_GE15","ITG1",2011,14.3,"Sicilia"
"Y_GE15","ITG2",2011,13.5,"Sardegna"
"Y_GE15","ITH",2011,5,"Nord-Est"
"Y_GE15","ITH1",2011,3.3,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2011,4.4,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2011,4.9,"Veneto"
"Y_GE15","ITH4",2011,5.2,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2011,5.2,"Emilia-Romagna"
"Y_GE15","ITI",2011,7.5,"Centro (IT)"
"Y_GE15","ITI1",2011,6.3,"Toscana"
"Y_GE15","ITI2",2011,6.4,"Umbria"
"Y_GE15","ITI3",2011,6.8,"Marche"
"Y_GE15","ITI4",2011,8.7,"Lazio"
"Y_GE15","LT",2011,15.4,"Lithuania"
"Y_GE15","LT0",2011,15.4,"Lietuva"
"Y_GE15","LT00",2011,15.4,"Lietuva"
"Y_GE15","LU",2011,4.9,"Luxembourg"
"Y_GE15","LU0",2011,4.9,"Luxembourg"
"Y_GE15","LU00",2011,4.9,"Luxembourg"
"Y_GE15","LV",2011,16.2,"Latvia"
"Y_GE15","LV0",2011,16.2,"Latvija"
"Y_GE15","LV00",2011,16.2,"Latvija"
"Y_GE15","MK",2011,31.4,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2011,31.4,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2011,31.4,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2011,6.4,"Malta"
"Y_GE15","MT0",2011,6.4,"Malta"
"Y_GE15","MT00",2011,6.4,"Malta"
"Y_GE15","NL",2011,5,"Netherlands"
"Y_GE15","NL1",2011,5.7,"Noord-Nederland"
"Y_GE15","NL11",2011,6.8,"Groningen"
"Y_GE15","NL12",2011,5.1,"Friesland (NL)"
"Y_GE15","NL13",2011,5.3,"Drenthe"
"Y_GE15","NL2",2011,4.8,"Oost-Nederland"
"Y_GE15","NL21",2011,4.9,"Overijssel"
"Y_GE15","NL22",2011,4.7,"Gelderland"
"Y_GE15","NL23",2011,5.4,"Flevoland"
"Y_GE15","NL3",2011,5,"West-Nederland"
"Y_GE15","NL31",2011,4.2,"Utrecht"
"Y_GE15","NL32",2011,5,"Noord-Holland"
"Y_GE15","NL33",2011,5.6,"Zuid-Holland"
"Y_GE15","NL34",2011,3.2,"Zeeland"
"Y_GE15","NL4",2011,4.7,"Zuid-Nederland"
"Y_GE15","NL41",2011,4.6,"Noord-Brabant"
"Y_GE15","NL42",2011,4.8,"Limburg (NL)"
"Y_GE15","NO",2011,3.2,"Norway"
"Y_GE15","NO0",2011,3.2,"Norge"
"Y_GE15","NO01",2011,3.4,"Oslo og Akershus"
"Y_GE15","NO02",2011,2.9,"Hedmark og Oppland"
"Y_GE15","NO03",2011,3.6,"Sør-Østlandet"
"Y_GE15","NO04",2011,2.2,"Agder og Rogaland"
"Y_GE15","NO05",2011,3.1,"Vestlandet"
"Y_GE15","NO06",2011,3.5,"Trøndelag"
"Y_GE15","NO07",2011,3.5,"Nord-Norge"
"Y_GE15","PL",2011,9.6,"Poland"
"Y_GE15","PL1",2011,8.3,"Region Centralny"
"Y_GE15","PL11",2011,9.3,"Lódzkie"
"Y_GE15","PL12",2011,7.9,"Mazowieckie"
"Y_GE15","PL2",2011,9.3,"Region Poludniowy"
"Y_GE15","PL21",2011,9.3,"Malopolskie"
"Y_GE15","PL22",2011,9.2,"Slaskie"
"Y_GE15","PL3",2011,11.3,"Region Wschodni"
"Y_GE15","PL31",2011,10.3,"Lubelskie"
"Y_GE15","PL32",2011,12.4,"Podkarpackie"
"Y_GE15","PL33",2011,12.9,"Swietokrzyskie"
"Y_GE15","PL34",2011,9.3,"Podlaskie"
"Y_GE15","PL4",2011,9.5,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2011,8.6,"Wielkopolskie"
"Y_GE15","PL42",2011,11.8,"Zachodniopomorskie"
"Y_GE15","PL43",2011,9.4,"Lubuskie"
"Y_GE15","PL5",2011,10.3,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2011,10.6,"Dolnoslaskie"
"Y_GE15","PL52",2011,9.3,"Opolskie"
"Y_GE15","PL6",2011,9.7,"Region Pólnocny"
"Y_GE15","PL61",2011,11,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2011,9.6,"Warminsko-Mazurskie"
"Y_GE15","PL63",2011,8.5,"Pomorskie"
"Y_GE15","PT",2011,12.7,"Portugal"
"Y_GE15","PT1",2011,12.7,"Continente"
"Y_GE15","PT11",2011,13,"Norte"
"Y_GE15","PT15",2011,15.4,"Algarve"
"Y_GE15","PT16",2011,10,"Centro (PT)"
"Y_GE15","PT17",2011,14.1,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2011,12.4,"Alentejo"
"Y_GE15","PT2",2011,11.3,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2011,11.3,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2011,13.5,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2011,13.5,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2011,7.2,"Romania"
"Y_GE15","RO1",2011,7.7,"Macroregiunea unu"
"Y_GE15","RO11",2011,5.1,"Nord-Vest"
"Y_GE15","RO12",2011,10.8,"Centru"
"Y_GE15","RO2",2011,6.7,"Macroregiunea doi"
"Y_GE15","RO21",2011,4.7,"Nord-Est"
"Y_GE15","RO22",2011,9.6,"Sud-Est"
"Y_GE15","RO3",2011,8,"Macroregiunea trei"
"Y_GE15","RO31",2011,10,"Sud - Muntenia"
"Y_GE15","RO32",2011,5.6,"Bucuresti - Ilfov"
"Y_GE15","RO4",2011,6.2,"Macroregiunea patru"
"Y_GE15","RO41",2011,6.6,"Sud-Vest Oltenia"
"Y_GE15","RO42",2011,5.7,"Vest"
"Y_GE15","SE",2011,7.8,"Sweden"
"Y_GE15","SE1",2011,7.3,"Östra Sverige"
"Y_GE15","SE11",2011,6.6,"Stockholm"
"Y_GE15","SE12",2011,8.4,"Östra Mellansverige"
"Y_GE15","SE2",2011,8,"Södra Sverige"
"Y_GE15","SE21",2011,7.1,"Småland med öarna"
"Y_GE15","SE22",2011,9.2,"Sydsverige"
"Y_GE15","SE23",2011,7.4,"Västsverige"
"Y_GE15","SE3",2011,8.5,"Norra Sverige"
"Y_GE15","SE31",2011,8.8,"Norra Mellansverige"
"Y_GE15","SE32",2011,8.8,"Mellersta Norrland"
"Y_GE15","SE33",2011,8,"Övre Norrland"
"Y_GE15","SI",2011,8.2,"Slovenia"
"Y_GE15","SI0",2011,8.2,"Slovenija"
"Y_GE15","SI03",2011,9.2,"Vzhodna Slovenija"
"Y_GE15","SI04",2011,7,"Zahodna Slovenija"
"Y_GE15","SK",2011,13.6,"Slovakia"
"Y_GE15","SK0",2011,13.6,"Slovensko"
"Y_GE15","SK01",2011,5.8,"Bratislavský kraj"
"Y_GE15","SK02",2011,10.7,"Západné Slovensko"
"Y_GE15","SK03",2011,15.9,"Stredné Slovensko"
"Y_GE15","SK04",2011,18.7,"Východné Slovensko"
"Y_GE15","TR",2011,8.8,"Turkey"
"Y_GE15","TR1",2011,11.1,"Istanbul"
"Y_GE15","TR10",2011,11.1,"Istanbul"
"Y_GE15","TR2",2011,6.3,"Bati Marmara"
"Y_GE15","TR21",2011,8.1,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2011,4.3,"Balikesir, Çanakkale"
"Y_GE15","TR3",2011,9.2,"Ege"
"Y_GE15","TR31",2011,13.7,"Izmir"
"Y_GE15","TR32",2011,7.5,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2011,4.5,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2011,8.7,"Dogu Marmara"
"Y_GE15","TR41",2011,6.7,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2011,10.6,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2011,7.5,"Bati Anadolu"
"Y_GE15","TR51",2011,8.5,"Ankara"
"Y_GE15","TR52",2011,5.5,"Konya, Karaman"
"Y_GE15","TR6",2011,9.4,"Akdeniz"
"Y_GE15","TR61",2011,8.7,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2011,9.3,"Adana, Mersin"
"Y_GE15","TR63",2011,10.5,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2011,8.7,"Orta Anadolu"
"Y_GE15","TR71",2011,7,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2011,9.8,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2011,5.3,"Bati Karadeniz"
"Y_GE15","TR81",2011,6.9,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2011,5.3,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2011,4.7,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2011,5.3,"Dogu Karadeniz"
"Y_GE15","TR90",2011,5.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2011,7.4,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2011,5.6,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2011,9.1,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2011,9.4,"Ortadogu Anadolu"
"Y_GE15","TRB1",2011,7.8,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2011,11,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2011,10.1,"Güneydogu Anadolu"
"Y_GE15","TRC1",2011,13.2,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2011,6.8,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2011,10.3,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2011,8,"United Kingdom"
"Y_GE15","UKC",2011,10.7,"North East (UK)"
"Y_GE15","UKC1",2011,11.8,"Tees Valley and Durham"
"Y_GE15","UKC2",2011,9.8,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2011,8.4,"North West (UK)"
"Y_GE15","UKD1",2011,7,"Cumbria"
"Y_GE15","UKD3",2011,9.7,"Greater Manchester"
"Y_GE15","UKD4",2011,6.8,"Lancashire"
"Y_GE15","UKD6",2011,5.7,"Cheshire"
"Y_GE15","UKD7",2011,10,"Merseyside"
"Y_GE15","UKE",2011,9.3,"Yorkshire and The Humber"
"Y_GE15","UKE1",2011,8.9,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2011,6.5,"North Yorkshire"
"Y_GE15","UKE3",2011,10.6,"South Yorkshire"
"Y_GE15","UKE4",2011,9.7,"West Yorkshire"
"Y_GE15","UKF",2011,7.9,"East Midlands (UK)"
"Y_GE15","UKF1",2011,8.8,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2011,7.5,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2011,6.5,"Lincolnshire"
"Y_GE15","UKG",2011,9,"West Midlands (UK)"
"Y_GE15","UKG1",2011,6.1,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2011,7.9,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2011,11.3,"West Midlands"
"Y_GE15","UKH",2011,6.6,"East of England"
"Y_GE15","UKH1",2011,6.3,"East Anglia"
"Y_GE15","UKH2",2011,6.7,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2011,6.8,"Essex"
"Y_GE15","UKI",2011,9.8,"London"
"Y_GE15","UKI3",2011,7.7,"Inner London - West"
"Y_GE15","UKI4",2011,12,"Inner London - East"
"Y_GE15","UKI5",2011,11.1,"Outer London - East and North East"
"Y_GE15","UKI6",2011,8.2,"Outer London - South"
"Y_GE15","UKI7",2011,8.5,"Outer London - West and North West"
"Y_GE15","UKJ",2011,6,"South East (UK)"
"Y_GE15","UKJ1",2011,5.2,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2011,5.3,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2011,6,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2011,8.2,"Kent"
"Y_GE15","UKK",2011,6.3,"South West (UK)"
"Y_GE15","UKK1",2011,6.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2011,6,"Dorset and Somerset"
"Y_GE15","UKK3",2011,6.2,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2011,6.5,"Devon"
"Y_GE15","UKL",2011,8.6,"Wales"
"Y_GE15","UKL1",2011,9.9,"West Wales and The Valleys"
"Y_GE15","UKL2",2011,6.5,"East Wales"
"Y_GE15","UKM",2011,8,"Scotland"
"Y_GE15","UKM2",2011,7.4,"Eastern Scotland"
"Y_GE15","UKM3",2011,9.6,"South Western Scotland"
"Y_GE15","UKM5",2011,4.6,"North Eastern Scotland"
"Y_GE15","UKM6",2011,6.9,"Highlands and Islands"
"Y_GE15","UKN",2011,7.2,"Northern Ireland (UK)"
"Y_GE15","UKN0",2011,7.2,"Northern Ireland (UK)"
"Y_GE25","AT",2011,3.9,"Austria"
"Y_GE25","AT1",2011,5.2,"Ostösterreich"
"Y_GE25","AT11",2011,3.3,"Burgenland (AT)"
"Y_GE25","AT12",2011,3.8,"Niederösterreich"
"Y_GE25","AT13",2011,6.8,"Wien"
"Y_GE25","AT2",2011,3.4,"Südösterreich"
"Y_GE25","AT21",2011,3.6,"Kärnten"
"Y_GE25","AT22",2011,3.4,"Steiermark"
"Y_GE25","AT3",2011,2.6,"Westösterreich"
"Y_GE25","AT31",2011,2.7,"Oberösterreich"
"Y_GE25","AT32",2011,2.4,"Salzburg"
"Y_GE25","AT33",2011,2.2,"Tirol"
"Y_GE25","AT34",2011,3.1,"Vorarlberg"
"Y_GE25","BE",2011,6,"Belgium"
"Y_GE25","BE1",2011,15.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2011,15.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2011,3.5,"Vlaams Gewest"
"Y_GE25","BE21",2011,4.7,"Prov. Antwerpen"
"Y_GE25","BE22",2011,3.7,"Prov. Limburg (BE)"
"Y_GE25","BE23",2011,3.1,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2011,2.9,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2011,2.4,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2011,7.9,"Région wallonne"
"Y_GE25","BE31",2011,5.6,"Prov. Brabant Wallon"
"Y_GE25","BE32",2011,9.6,"Prov. Hainaut"
"Y_GE25","BE33",2011,8,"Prov. Liège"
"Y_GE25","BE34",2011,4.9,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2011,6.5,"Prov. Namur"
"Y_GE25","BG",2011,10.1,"Bulgaria"
"Y_GE25","BG3",2011,11.8,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2011,11.3,"Severozapaden"
"Y_GE25","BG32",2011,11.4,"Severen tsentralen"
"Y_GE25","BG33",2011,14.2,"Severoiztochen"
"Y_GE25","BG34",2011,10.3,"Yugoiztochen"
"Y_GE25","BG4",2011,8.5,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2011,6.7,"Yugozapaden"
"Y_GE25","BG42",2011,11.6,"Yuzhen tsentralen"
"Y_GE25","CH",2011,3.5,"Switzerland"
"Y_GE25","CH0",2011,3.5,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2011,5.1,"Région lémanique"
"Y_GE25","CH02",2011,2.9,"Espace Mittelland"
"Y_GE25","CH03",2011,3.6,"Nordwestschweiz"
"Y_GE25","CH04",2011,3.5,"Zürich"
"Y_GE25","CH05",2011,2.6,"Ostschweiz"
"Y_GE25","CH06",2011,2.1,"Zentralschweiz"
"Y_GE25","CH07",2011,4.5,"Ticino"
"Y_GE25","CY",2011,6.4,"Cyprus"
"Y_GE25","CY0",2011,6.4,"Kypros"
"Y_GE25","CY00",2011,6.4,"Kypros"
"Y_GE25","CZ",2011,5.8,"Czech Republic"
"Y_GE25","CZ0",2011,5.8,"Ceská republika"
"Y_GE25","CZ01",2011,3.2,"Praha"
"Y_GE25","CZ02",2011,4.2,"Strední Cechy"
"Y_GE25","CZ03",2011,4.6,"Jihozápad"
"Y_GE25","CZ04",2011,7.9,"Severozápad"
"Y_GE25","CZ05",2011,5.7,"Severovýchod"
"Y_GE25","CZ06",2011,6.3,"Jihovýchod"
"Y_GE25","CZ07",2011,6.7,"Strední Morava"
"Y_GE25","CZ08",2011,8.6,"Moravskoslezsko"
"Y_GE25","DE",2011,5.5,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2011,3.3,"Baden-Württemberg"
"Y_GE25","DE11",2011,3.3,"Stuttgart"
"Y_GE25","DE12",2011,3.9,"Karlsruhe"
"Y_GE25","DE13",2011,2.7,"Freiburg"
"Y_GE25","DE14",2011,2.9,"Tübingen"
"Y_GE25","DE2",2011,3,"Bayern"
"Y_GE25","DE21",2011,2.5,"Oberbayern"
"Y_GE25","DE22",2011,2.4,"Niederbayern"
"Y_GE25","DE23",2011,3.1,"Oberpfalz"
"Y_GE25","DE24",2011,3.8,"Oberfranken"
"Y_GE25","DE25",2011,3.7,"Mittelfranken"
"Y_GE25","DE26",2011,3.3,"Unterfranken"
"Y_GE25","DE27",2011,2.9,"Schwaben"
"Y_GE25","DE3",2011,11.5,"Berlin"
"Y_GE25","DE30",2011,11.5,"Berlin"
"Y_GE25","DE4",2011,8.4,"Brandenburg"
"Y_GE25","DE40",2011,8.4,"Brandenburg"
"Y_GE25","DE5",2011,6.8,"Bremen"
"Y_GE25","DE50",2011,6.8,"Bremen"
"Y_GE25","DE6",2011,5.2,"Hamburg"
"Y_GE25","DE60",2011,5.2,"Hamburg"
"Y_GE25","DE7",2011,4.2,"Hessen"
"Y_GE25","DE71",2011,4.2,"Darmstadt"
"Y_GE25","DE72",2011,4.4,"Gießen"
"Y_GE25","DE73",2011,4.2,"Kassel"
"Y_GE25","DE8",2011,10,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2011,10,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2011,5,"Niedersachsen"
"Y_GE25","DE91",2011,5.6,"Braunschweig"
"Y_GE25","DE92",2011,6,"Hannover"
"Y_GE25","DE93",2011,4.8,"Lüneburg"
"Y_GE25","DE94",2011,3.9,"Weser-Ems"
"Y_GE25","DEA",2011,5.9,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2011,6.2,"Düsseldorf"
"Y_GE25","DEA2",2011,5.5,"Köln"
"Y_GE25","DEA3",2011,5.1,"Münster"
"Y_GE25","DEA4",2011,5,"Detmold"
"Y_GE25","DEA5",2011,6.8,"Arnsberg"
"Y_GE25","DEB",2011,4.2,"Rheinland-Pfalz"
"Y_GE25","DEB1",2011,4,"Koblenz"
"Y_GE25","DEB2",2011,3.3,"Trier"
"Y_GE25","DEB3",2011,4.5,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2011,5.3,"Saarland"
"Y_GE25","DEC0",2011,5.3,"Saarland"
"Y_GE25","DED",2011,9.2,"Sachsen"
"Y_GE25","DED2",2011,8.5,"Dresden"
"Y_GE25","DED4",2011,8.7,"Chemnitz"
"Y_GE25","DED5",2011,11,"Leipzig"
"Y_GE25","DEE",2011,10,"Sachsen-Anhalt"
"Y_GE25","DEE0",2011,10,"Sachsen-Anhalt"
"Y_GE25","DEF",2011,5.4,"Schleswig-Holstein"
"Y_GE25","DEF0",2011,5.4,"Schleswig-Holstein"
"Y_GE25","DEG",2011,7.5,"Thüringen"
"Y_GE25","DEG0",2011,7.5,"Thüringen"
"Y_GE25","DK",2011,6.3,"Denmark"
"Y_GE25","DK0",2011,6.3,"Danmark"
"Y_GE25","DK01",2011,6.8,"Hovedstaden"
"Y_GE25","DK02",2011,5.9,"Sjælland"
"Y_GE25","DK03",2011,6.4,"Syddanmark"
"Y_GE25","DK04",2011,5.6,"Midtjylland"
"Y_GE25","DK05",2011,6.8,"Nordjylland"
"Y_GE25","EA17",2011,8.9,"Euro area (17 countries)"
"Y_GE25","EA18",2011,8.9,"Euro area (18 countries)"
"Y_GE25","EA19",2011,9,"Euro area (19 countries)"
"Y_GE25","EE",2011,11.2,"Estonia"
"Y_GE25","EE0",2011,11.2,"Eesti"
"Y_GE25","EE00",2011,11.2,"Eesti"
"Y_GE25","EL",2011,15.9,"Greece"
"Y_GE25","EL3",2011,16.3,"Attiki"
"Y_GE25","EL30",2011,16.3,"Attiki"
"Y_GE25","EL4",2011,13.4,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2011,12.6,"Voreio Aigaio"
"Y_GE25","EL42",2011,13.2,"Notio Aigaio"
"Y_GE25","EL43",2011,13.6,"Kriti"
"Y_GE25","EL5",2011,17.6,"Voreia Ellada"
"Y_GE25","EL51",2011,17.2,"Anatoliki Makedonia, Thraki"
"Y_GE25","EL52",2011,17.8,"Kentriki Makedonia"
"Y_GE25","EL53",2011,21.1,"Dytiki Makedonia"
"Y_GE25","EL54",2011,14.2,"Ipeiros"
"Y_GE25","EL6",2011,14.5,"Kentriki Ellada"
"Y_GE25","EL61",2011,14.4,"Thessalia"
"Y_GE25","EL62",2011,13.4,"Ionia Nisia"
"Y_GE25","EL63",2011,14.9,"Dytiki Ellada"
"Y_GE25","EL64",2011,16.9,"Sterea Ellada"
"Y_GE25","EL65",2011,12.4,"Peloponnisos"
"Y_GE25","ES",2011,19.2,"Spain"
"Y_GE25","ES1",2011,15.6,"Noroeste (ES)"
"Y_GE25","ES11",2011,15.8,"Galicia"
"Y_GE25","ES12",2011,16,"Principado de Asturias"
"Y_GE25","ES13",2011,13.6,"Cantabria"
"Y_GE25","ES2",2011,12.6,"Noreste (ES)"
"Y_GE25","ES21",2011,10.9,"País Vasco"
"Y_GE25","ES22",2011,11.7,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2011,14.9,"La Rioja"
"Y_GE25","ES24",2011,15.3,"Aragón"
"Y_GE25","ES3",2011,14.4,"Comunidad de Madrid"
"Y_GE25","ES30",2011,14.4,"Comunidad de Madrid"
"Y_GE25","ES4",2011,18.4,"Centro (ES)"
"Y_GE25","ES41",2011,15.1,"Castilla y León"
"Y_GE25","ES42",2011,20.4,"Castilla-la Mancha"
"Y_GE25","ES43",2011,22.2,"Extremadura"
"Y_GE25","ES5",2011,18.8,"Este (ES)"
"Y_GE25","ES51",2011,16.9,"Cataluña"
"Y_GE25","ES52",2011,21.5,"Comunidad Valenciana"
"Y_GE25","ES53",2011,19.9,"Illes Balears"
"Y_GE25","ES6",2011,26.6,"Sur (ES)"
"Y_GE25","ES61",2011,27.5,"Andalucía"
"Y_GE25","ES62",2011,22.5,"Región de Murcia"
"Y_GE25","ES63",2011,22.8,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2011,19,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2011,27.3,"Canarias (ES)"
"Y_GE25","ES70",2011,27.3,"Canarias (ES)"
"Y_GE25","EU15",2011,8.3,"European Union (15 countries)"
"Y_GE25","EU27",2011,8.2,"European Union (27 countries)"
"Y_GE25","EU28",2011,8.3,"European Union (28 countries)"
"Y_GE25","FI",2011,6.1,"Finland"
"Y_GE25","FI1",2011,6.1,"Manner-Suomi"
"Y_GE25","FI19",2011,6.2,"Länsi-Suomi"
"Y_GE25","FI1B",2011,4.7,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2011,6.9,"Etelä-Suomi"
"Y_GE25","FI1D",2011,7.4,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2011,NA,"Åland"
"Y_GE25","FI20",2011,NA,"Åland"
"Y_GE25","FR",2011,7.7,"France"
"Y_GE25","FR1",2011,7.3,"Île de France"
"Y_GE25","FR10",2011,7.3,"Île de France"
"Y_GE25","FR2",2011,7.2,"Bassin Parisien"
"Y_GE25","FR21",2011,8.2,"Champagne-Ardenne"
"Y_GE25","FR22",2011,7.3,"Picardie"
"Y_GE25","FR23",2011,7.2,"Haute-Normandie"
"Y_GE25","FR24",2011,6.9,"Centre (FR)"
"Y_GE25","FR25",2011,7.2,"Basse-Normandie"
"Y_GE25","FR26",2011,7,"Bourgogne"
"Y_GE25","FR3",2011,9.9,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2011,9.9,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2011,7.2,"Est (FR)"
"Y_GE25","FR41",2011,8.8,"Lorraine"
"Y_GE25","FR42",2011,5.7,"Alsace"
"Y_GE25","FR43",2011,6.8,"Franche-Comté"
"Y_GE25","FR5",2011,6.7,"Ouest (FR)"
"Y_GE25","FR51",2011,7.3,"Pays de la Loire"
"Y_GE25","FR52",2011,5.9,"Bretagne"
"Y_GE25","FR53",2011,6.7,"Poitou-Charentes"
"Y_GE25","FR6",2011,7,"Sud-Ouest (FR)"
"Y_GE25","FR61",2011,7.5,"Aquitaine"
"Y_GE25","FR62",2011,6.7,"Midi-Pyrénées"
"Y_GE25","FR63",2011,6.1,"Limousin"
"Y_GE25","FR7",2011,6.4,"Centre-Est (FR)"
"Y_GE25","FR71",2011,6.3,"Rhône-Alpes"
"Y_GE25","FR72",2011,6.6,"Auvergne"
"Y_GE25","FR8",2011,8.8,"Méditerranée"
"Y_GE25","FR81",2011,9.9,"Languedoc-Roussillon"
"Y_GE25","FR82",2011,8.4,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2011,NA,"Corse"
"Y_GE25","FRA",2011,21.6,"Départements d'outre-mer"
"Y_GE25","FRA1",2011,20.2,"Guadeloupe"
"Y_GE25","FRA2",2011,17.5,"Martinique"
"Y_GE25","FRA3",2011,18.1,"Guyane"
"Y_GE25","FRA4",2011,25.2,"La Réunion"
"Y_GE25","HR",2011,11.5,"Croatia"
"Y_GE25","HR0",2011,11.5,"Hrvatska"
"Y_GE25","HR03",2011,11.5,"Jadranska Hrvatska"
"Y_GE25","HR04",2011,11.5,"Kontinentalna Hrvatska"
"Y_GE25","HU",2011,9.9,"Hungary"
"Y_GE25","HU1",2011,8.3,"Közép-Magyarország"
"Y_GE25","HU10",2011,8.3,"Közép-Magyarország"
"Y_GE25","HU2",2011,8.8,"Dunántúl"
"Y_GE25","HU21",2011,8.5,"Közép-Dunántúl"
"Y_GE25","HU22",2011,6.6,"Nyugat-Dunántúl"
"Y_GE25","HU23",2011,11.8,"Dél-Dunántúl"
"Y_GE25","HU3",2011,12.2,"Alföld és Észak"
"Y_GE25","HU31",2011,14.8,"Észak-Magyarország"
"Y_GE25","HU32",2011,12.9,"Észak-Alföld"
"Y_GE25","HU33",2011,9.3,"Dél-Alföld"
"Y_GE25","IE",2011,12.8,"Ireland"
"Y_GE25","IE0",2011,12.8,"Éire/Ireland"
"Y_GE25","IE01",2011,13.8,"Border, Midland and Western"
"Y_GE25","IE02",2011,12.5,"Southern and Eastern"
"Y_GE25","IS",2011,5.5,"Iceland"
"Y_GE25","IS0",2011,5.5,"Ísland"
"Y_GE25","IS00",2011,5.5,"Ísland"
"Y_GE25","IT",2011,6.9,"Italy"
"Y_GE25","ITC",2011,5.2,"Nord-Ovest"
"Y_GE25","ITC1",2011,6.4,"Piemonte"
"Y_GE25","ITC2",2011,4.3,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2011,5.3,"Liguria"
"Y_GE25","ITC4",2011,4.7,"Lombardia"
"Y_GE25","ITF",2011,11.1,"Sud"
"Y_GE25","ITF1",2011,7.4,"Abruzzo"
"Y_GE25","ITF2",2011,8.6,"Molise"
"Y_GE25","ITF3",2011,12.9,"Campania"
"Y_GE25","ITF4",2011,10.8,"Puglia"
"Y_GE25","ITF5",2011,9.9,"Basilicata"
"Y_GE25","ITF6",2011,10.6,"Calabria"
"Y_GE25","ITG",2011,11.6,"Isole"
"Y_GE25","ITG1",2011,11.7,"Sicilia"
"Y_GE25","ITG2",2011,11.3,"Sardegna"
"Y_GE25","ITH",2011,4,"Nord-Est"
"Y_GE25","ITH1",2011,2.7,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2011,3.7,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2011,3.8,"Veneto"
"Y_GE25","ITH4",2011,4.2,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2011,4.3,"Emilia-Romagna"
"Y_GE25","ITI",2011,6.2,"Centro (IT)"
"Y_GE25","ITI1",2011,5.3,"Toscana"
"Y_GE25","ITI2",2011,5.3,"Umbria"
"Y_GE25","ITI3",2011,5.8,"Marche"
"Y_GE25","ITI4",2011,7.1,"Lazio"
"Y_GE25","LT",2011,13.9,"Lithuania"
"Y_GE25","LT0",2011,13.9,"Lietuva"
"Y_GE25","LT00",2011,13.9,"Lietuva"
"Y_GE25","LU",2011,4.1,"Luxembourg"
"Y_GE25","LU0",2011,4.1,"Luxembourg"
"Y_GE25","LU00",2011,4.1,"Luxembourg"
"Y_GE25","LV",2011,14.6,"Latvia"
"Y_GE25","LV0",2011,14.6,"Latvija"
"Y_GE25","LV00",2011,14.6,"Latvija"
"Y_GE25","MK",2011,28.5,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2011,28.5,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2011,28.5,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2011,5,"Malta"
"Y_GE25","MT0",2011,5,"Malta"
"Y_GE25","MT00",2011,5,"Malta"
"Y_GE25","NL",2011,4,"Netherlands"
"Y_GE25","NL1",2011,4.5,"Noord-Nederland"
"Y_GE25","NL11",2011,5.4,"Groningen"
"Y_GE25","NL12",2011,4.1,"Friesland (NL)"
"Y_GE25","NL13",2011,4.2,"Drenthe"
"Y_GE25","NL2",2011,3.9,"Oost-Nederland"
"Y_GE25","NL21",2011,3.8,"Overijssel"
"Y_GE25","NL22",2011,3.9,"Gelderland"
"Y_GE25","NL23",2011,4.7,"Flevoland"
"Y_GE25","NL3",2011,4.1,"West-Nederland"
"Y_GE25","NL31",2011,3.5,"Utrecht"
"Y_GE25","NL32",2011,4,"Noord-Holland"
"Y_GE25","NL33",2011,4.6,"Zuid-Holland"
"Y_GE25","NL34",2011,2.7,"Zeeland"
"Y_GE25","NL4",2011,3.8,"Zuid-Nederland"
"Y_GE25","NL41",2011,3.7,"Noord-Brabant"
"Y_GE25","NL42",2011,3.9,"Limburg (NL)"
"Y_GE25","NO",2011,2.4,"Norway"
"Y_GE25","NO0",2011,2.4,"Norge"
"Y_GE25","NO01",2011,2.6,"Oslo og Akershus"
"Y_GE25","NO02",2011,2.4,"Hedmark og Oppland"
"Y_GE25","NO03",2011,2.7,"Sør-Østlandet"
"Y_GE25","NO04",2011,1.5,"Agder og Rogaland"
"Y_GE25","NO05",2011,2.3,"Vestlandet"
"Y_GE25","NO06",2011,2.5,"Trøndelag"
"Y_GE25","NO07",2011,2.4,"Nord-Norge"
"Y_GE25","PL",2011,8,"Poland"
"Y_GE25","PL1",2011,6.9,"Region Centralny"
"Y_GE25","PL11",2011,7.9,"Lódzkie"
"Y_GE25","PL12",2011,6.4,"Mazowieckie"
"Y_GE25","PL2",2011,7.7,"Region Poludniowy"
"Y_GE25","PL21",2011,7.8,"Malopolskie"
"Y_GE25","PL22",2011,7.7,"Slaskie"
"Y_GE25","PL3",2011,9.1,"Region Wschodni"
"Y_GE25","PL31",2011,8.1,"Lubelskie"
"Y_GE25","PL32",2011,10,"Podkarpackie"
"Y_GE25","PL33",2011,10.6,"Swietokrzyskie"
"Y_GE25","PL34",2011,7.6,"Podlaskie"
"Y_GE25","PL4",2011,7.7,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2011,6.8,"Wielkopolskie"
"Y_GE25","PL42",2011,9.8,"Zachodniopomorskie"
"Y_GE25","PL43",2011,8,"Lubuskie"
"Y_GE25","PL5",2011,8.9,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2011,9.2,"Dolnoslaskie"
"Y_GE25","PL52",2011,8,"Opolskie"
"Y_GE25","PL6",2011,8,"Region Pólnocny"
"Y_GE25","PL61",2011,9.2,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2011,7.9,"Warminsko-Mazurskie"
"Y_GE25","PL63",2011,7,"Pomorskie"
"Y_GE25","PT",2011,11.1,"Portugal"
"Y_GE25","PT1",2011,11.2,"Continente"
"Y_GE25","PT11",2011,11.5,"Norte"
"Y_GE25","PT15",2011,13.7,"Algarve"
"Y_GE25","PT16",2011,8.8,"Centro (PT)"
"Y_GE25","PT17",2011,12.5,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2011,10.9,"Alentejo"
"Y_GE25","PT2",2011,8.7,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2011,8.7,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2011,11.1,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2011,11.1,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2011,5.7,"Romania"
"Y_GE25","RO1",2011,5.8,"Macroregiunea unu"
"Y_GE25","RO11",2011,3.7,"Nord-Vest"
"Y_GE25","RO12",2011,8.5,"Centru"
"Y_GE25","RO2",2011,5.5,"Macroregiunea doi"
"Y_GE25","RO21",2011,3.9,"Nord-Est"
"Y_GE25","RO22",2011,7.8,"Sud-Est"
"Y_GE25","RO3",2011,6.1,"Macroregiunea trei"
"Y_GE25","RO31",2011,7.7,"Sud - Muntenia"
"Y_GE25","RO32",2011,4.3,"Bucuresti - Ilfov"
"Y_GE25","RO4",2011,5.1,"Macroregiunea patru"
"Y_GE25","RO41",2011,5.6,"Sud-Vest Oltenia"
"Y_GE25","RO42",2011,4.4,"Vest"
"Y_GE25","SE",2011,5.5,"Sweden"
"Y_GE25","SE1",2011,5.3,"Östra Sverige"
"Y_GE25","SE11",2011,4.8,"Stockholm"
"Y_GE25","SE12",2011,6,"Östra Mellansverige"
"Y_GE25","SE2",2011,5.7,"Södra Sverige"
"Y_GE25","SE21",2011,4.9,"Småland med öarna"
"Y_GE25","SE22",2011,6.8,"Sydsverige"
"Y_GE25","SE23",2011,5.2,"Västsverige"
"Y_GE25","SE3",2011,5.8,"Norra Sverige"
"Y_GE25","SE31",2011,6.2,"Norra Mellansverige"
"Y_GE25","SE32",2011,5.5,"Mellersta Norrland"
"Y_GE25","SE33",2011,5.2,"Övre Norrland"
"Y_GE25","SI",2011,7.5,"Slovenia"
"Y_GE25","SI0",2011,7.5,"Slovenija"
"Y_GE25","SI03",2011,8.4,"Vzhodna Slovenija"
"Y_GE25","SI04",2011,6.4,"Zahodna Slovenija"
"Y_GE25","SK",2011,11.8,"Slovakia"
"Y_GE25","SK0",2011,11.8,"Slovensko"
"Y_GE25","SK01",2011,5.1,"Bratislavský kraj"
"Y_GE25","SK02",2011,9.3,"Západné Slovensko"
"Y_GE25","SK03",2011,13.7,"Stredné Slovensko"
"Y_GE25","SK04",2011,16.2,"Východné Slovensko"
"Y_GE25","TR",2011,7.2,"Turkey"
"Y_GE25","TR1",2011,9.6,"Istanbul"
"Y_GE25","TR10",2011,9.6,"Istanbul"
"Y_GE25","TR2",2011,4.9,"Bati Marmara"
"Y_GE25","TR21",2011,6.4,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2011,3.3,"Balikesir, Çanakkale"
"Y_GE25","TR3",2011,7.4,"Ege"
"Y_GE25","TR31",2011,11.3,"Izmir"
"Y_GE25","TR32",2011,5.9,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2011,3.3,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2011,7.2,"Dogu Marmara"
"Y_GE25","TR41",2011,5.5,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2011,8.9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2011,6,"Bati Anadolu"
"Y_GE25","TR51",2011,6.7,"Ankara"
"Y_GE25","TR52",2011,4.3,"Konya, Karaman"
"Y_GE25","TR6",2011,7.9,"Akdeniz"
"Y_GE25","TR61",2011,7.3,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2011,7.7,"Adana, Mersin"
"Y_GE25","TR63",2011,8.9,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2011,7,"Orta Anadolu"
"Y_GE25","TR71",2011,5.5,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2011,7.9,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2011,4.2,"Bati Karadeniz"
"Y_GE25","TR81",2011,4.8,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2011,4.4,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2011,3.8,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2011,3.6,"Dogu Karadeniz"
"Y_GE25","TR90",2011,3.6,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2011,6.1,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2011,4.2,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2011,7.8,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2011,7.7,"Ortadogu Anadolu"
"Y_GE25","TRB1",2011,5.8,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2011,9.7,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2011,8.6,"Güneydogu Anadolu"
"Y_GE25","TRC1",2011,11.1,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2011,6.1,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2011,8.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2011,5.8,"United Kingdom"
"Y_GE25","UKC",2011,8.5,"North East (UK)"
"Y_GE25","UKC1",2011,9.6,"Tees Valley and Durham"
"Y_GE25","UKC2",2011,7.6,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2011,5.6,"North West (UK)"
"Y_GE25","UKD1",2011,4.3,"Cumbria"
"Y_GE25","UKD3",2011,6.6,"Greater Manchester"
"Y_GE25","UKD4",2011,4,"Lancashire"
"Y_GE25","UKD6",2011,3.9,"Cheshire"
"Y_GE25","UKD7",2011,6.9,"Merseyside"
"Y_GE25","UKE",2011,6.7,"Yorkshire and The Humber"
"Y_GE25","UKE1",2011,6.6,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2011,4.4,"North Yorkshire"
"Y_GE25","UKE3",2011,7.2,"South Yorkshire"
"Y_GE25","UKE4",2011,7.3,"West Yorkshire"
"Y_GE25","UKF",2011,5.6,"East Midlands (UK)"
"Y_GE25","UKF1",2011,6.1,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2011,5.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2011,4.8,"Lincolnshire"
"Y_GE25","UKG",2011,6.4,"West Midlands (UK)"
"Y_GE25","UKG1",2011,4.1,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2011,5.8,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2011,8.1,"West Midlands"
"Y_GE25","UKH",2011,4.8,"East of England"
"Y_GE25","UKH1",2011,4.6,"East Anglia"
"Y_GE25","UKH2",2011,5.2,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2011,4.5,"Essex"
"Y_GE25","UKI",2011,7.8,"London"
"Y_GE25","UKI3",2011,5.7,"Inner London - West"
"Y_GE25","UKI4",2011,9.4,"Inner London - East"
"Y_GE25","UKI5",2011,8.8,"Outer London - East and North East"
"Y_GE25","UKI6",2011,6.6,"Outer London - South"
"Y_GE25","UKI7",2011,7.2,"Outer London - West and North West"
"Y_GE25","UKJ",2011,4.3,"South East (UK)"
"Y_GE25","UKJ1",2011,4.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2011,3.9,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2011,4.3,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2011,5.6,"Kent"
"Y_GE25","UKK",2011,4.6,"South West (UK)"
"Y_GE25","UKK1",2011,4.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2011,4.6,"Dorset and Somerset"
"Y_GE25","UKK3",2011,5.4,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2011,4.4,"Devon"
"Y_GE25","UKL",2011,5.7,"Wales"
"Y_GE25","UKL1",2011,6.8,"West Wales and The Valleys"
"Y_GE25","UKL2",2011,3.9,"East Wales"
"Y_GE25","UKM",2011,5.4,"Scotland"
"Y_GE25","UKM2",2011,4.9,"Eastern Scotland"
"Y_GE25","UKM3",2011,6.5,"South Western Scotland"
"Y_GE25","UKM5",2011,3.1,"North Eastern Scotland"
"Y_GE25","UKM6",2011,5.7,"Highlands and Islands"
"Y_GE25","UKN",2011,5.2,"Northern Ireland (UK)"
"Y_GE25","UKN0",2011,5.2,"Northern Ireland (UK)"
"Y15-24","AT",2010,9.5,"Austria"
"Y15-24","AT1",2010,12.5,"Ostösterreich"
"Y15-24","AT11",2010,NA,"Burgenland (AT)"
"Y15-24","AT12",2010,7.4,"Niederösterreich"
"Y15-24","AT13",2010,18.1,"Wien"
"Y15-24","AT2",2010,8.8,"Südösterreich"
"Y15-24","AT21",2010,NA,"Kärnten"
"Y15-24","AT22",2010,9.1,"Steiermark"
"Y15-24","AT3",2010,7.2,"Westösterreich"
"Y15-24","AT31",2010,6.9,"Oberösterreich"
"Y15-24","AT32",2010,NA,"Salzburg"
"Y15-24","AT33",2010,6.6,"Tirol"
"Y15-24","AT34",2010,NA,"Vorarlberg"
"Y15-24","BE",2010,22.4,"Belgium"
"Y15-24","BE1",2010,39.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2010,39.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2010,15.6,"Vlaams Gewest"
"Y15-24","BE21",2010,18.2,"Prov. Antwerpen"
"Y15-24","BE22",2010,17.4,"Prov. Limburg (BE)"
"Y15-24","BE23",2010,15.7,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2010,15.1,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2010,11,"Prov. West-Vlaanderen"
"Y15-24","BE3",2010,30,"Région wallonne"
"Y15-24","BE31",2010,27.1,"Prov. Brabant Wallon"
"Y15-24","BE32",2010,35.9,"Prov. Hainaut"
"Y15-24","BE33",2010,27.3,"Prov. Liège"
"Y15-24","BE34",2010,19.9,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2010,28,"Prov. Namur"
"Y15-24","BG",2010,21.9,"Bulgaria"
"Y15-24","BG3",2010,24.3,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2010,22,"Severozapaden"
"Y15-24","BG32",2010,25.5,"Severen tsentralen"
"Y15-24","BG33",2010,24.7,"Severoiztochen"
"Y15-24","BG34",2010,24.6,"Yugoiztochen"
"Y15-24","BG4",2010,20.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2010,14.7,"Yugozapaden"
"Y15-24","BG42",2010,31.6,"Yuzhen tsentralen"
"Y15-24","CH",2010,7.9,"Switzerland"
"Y15-24","CH0",2010,7.9,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2010,12.9,"Région lémanique"
"Y15-24","CH02",2010,7.7,"Espace Mittelland"
"Y15-24","CH03",2010,8.1,"Nordwestschweiz"
"Y15-24","CH04",2010,6.8,"Zürich"
"Y15-24","CH05",2010,5.2,"Ostschweiz"
"Y15-24","CH06",2010,4.8,"Zentralschweiz"
"Y15-24","CH07",2010,10.7,"Ticino"
"Y15-24","CY",2010,16.6,"Cyprus"
"Y15-24","CY0",2010,16.6,"Kypros"
"Y15-24","CY00",2010,16.6,"Kypros"
"Y15-24","CZ",2010,18.3,"Czech Republic"
"Y15-24","CZ0",2010,18.3,"Ceská republika"
"Y15-24","CZ01",2010,8.8,"Praha"
"Y15-24","CZ02",2010,16,"Strední Cechy"
"Y15-24","CZ03",2010,15.6,"Jihozápad"
"Y15-24","CZ04",2010,26.4,"Severozápad"
"Y15-24","CZ05",2010,20.8,"Severovýchod"
"Y15-24","CZ06",2010,16.6,"Jihovýchod"
"Y15-24","CZ07",2010,19.9,"Strední Morava"
"Y15-24","CZ08",2010,20,"Moravskoslezsko"
"Y15-24","DE",2010,9.8,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2010,7,"Baden-Württemberg"
"Y15-24","DE11",2010,7.1,"Stuttgart"
"Y15-24","DE12",2010,8.8,"Karlsruhe"
"Y15-24","DE13",2010,5.4,"Freiburg"
"Y15-24","DE14",2010,6.2,"Tübingen"
"Y15-24","DE2",2010,6.5,"Bayern"
"Y15-24","DE21",2010,5,"Oberbayern"
"Y15-24","DE22",2010,6.4,"Niederbayern"
"Y15-24","DE23",2010,NA,"Oberpfalz"
"Y15-24","DE24",2010,9.2,"Oberfranken"
"Y15-24","DE25",2010,8.7,"Mittelfranken"
"Y15-24","DE26",2010,8.4,"Unterfranken"
"Y15-24","DE27",2010,5.5,"Schwaben"
"Y15-24","DE3",2010,16.5,"Berlin"
"Y15-24","DE30",2010,16.5,"Berlin"
"Y15-24","DE4",2010,14.7,"Brandenburg"
"Y15-24","DE40",2010,14.7,"Brandenburg"
"Y15-24","DE5",2010,NA,"Bremen"
"Y15-24","DE50",2010,NA,"Bremen"
"Y15-24","DE6",2010,7.3,"Hamburg"
"Y15-24","DE60",2010,7.3,"Hamburg"
"Y15-24","DE7",2010,11.1,"Hessen"
"Y15-24","DE71",2010,10.6,"Darmstadt"
"Y15-24","DE72",2010,13,"Gießen"
"Y15-24","DE73",2010,11,"Kassel"
"Y15-24","DE8",2010,13.3,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2010,13.3,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2010,10.4,"Niedersachsen"
"Y15-24","DE91",2010,10.4,"Braunschweig"
"Y15-24","DE92",2010,11.5,"Hannover"
"Y15-24","DE93",2010,10.9,"Lüneburg"
"Y15-24","DE94",2010,9.3,"Weser-Ems"
"Y15-24","DEA",2010,10.8,"Nordrhein-Westfalen"
"Y15-24","DEA1",2010,11.7,"Düsseldorf"
"Y15-24","DEA2",2010,10.4,"Köln"
"Y15-24","DEA3",2010,9.1,"Münster"
"Y15-24","DEA4",2010,10.5,"Detmold"
"Y15-24","DEA5",2010,11.7,"Arnsberg"
"Y15-24","DEB",2010,9.4,"Rheinland-Pfalz"
"Y15-24","DEB1",2010,6.6,"Koblenz"
"Y15-24","DEB2",2010,NA,"Trier"
"Y15-24","DEB3",2010,12.5,"Rheinhessen-Pfalz"
"Y15-24","DEC",2010,NA,"Saarland"
"Y15-24","DEC0",2010,NA,"Saarland"
"Y15-24","DED",2010,12.6,"Sachsen"
"Y15-24","DED2",2010,12.1,"Dresden"
"Y15-24","DED4",2010,11.8,"Chemnitz"
"Y15-24","DED5",2010,14.4,"Leipzig"
"Y15-24","DEE",2010,13.2,"Sachsen-Anhalt"
"Y15-24","DEE0",2010,13.2,"Sachsen-Anhalt"
"Y15-24","DEF",2010,10.2,"Schleswig-Holstein"
"Y15-24","DEF0",2010,10.2,"Schleswig-Holstein"
"Y15-24","DEG",2010,10.5,"Thüringen"
"Y15-24","DEG0",2010,10.5,"Thüringen"
"Y15-24","DK",2010,14,"Denmark"
"Y15-24","DK0",2010,14,"Danmark"
"Y15-24","DK01",2010,14.7,"Hovedstaden"
"Y15-24","DK02",2010,15.7,"Sjælland"
"Y15-24","DK03",2010,13.8,"Syddanmark"
"Y15-24","DK04",2010,13.4,"Midtjylland"
"Y15-24","DK05",2010,11.3,"Nordjylland"
"Y15-24","EA17",2010,20.8,"Euro area (17 countries)"
"Y15-24","EA18",2010,21,"Euro area (18 countries)"
"Y15-24","EA19",2010,21.1,"Euro area (19 countries)"
"Y15-24","EE",2010,32.9,"Estonia"
"Y15-24","EE0",2010,32.9,"Eesti"
"Y15-24","EE00",2010,32.9,"Eesti"
"Y15-24","EL",2010,33,"Greece"
"Y15-24","EL3",2010,30.9,"Attiki"
"Y15-24","EL30",2010,30.9,"Attiki"
"Y15-24","EL4",2010,29.6,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2010,29.7,"Voreio Aigaio"
"Y15-24","EL42",2010,28.4,"Notio Aigaio"
"Y15-24","EL43",2010,30.4,"Kriti"
"Y15-24","EL5",2010,36,"Voreia Ellada"
"Y15-24","EL51",2010,40.1,"Anatoliki Makedonia, Thraki"
"Y15-24","EL52",2010,34.1,"Kentriki Makedonia"
"Y15-24","EL53",2010,35.3,"Dytiki Makedonia"
"Y15-24","EL54",2010,37.1,"Ipeiros"
"Y15-24","EL6",2010,34.3,"Kentriki Ellada"
"Y15-24","EL61",2010,34.4,"Thessalia"
"Y15-24","EL62",2010,35.2,"Ionia Nisia"
"Y15-24","EL63",2010,35.3,"Dytiki Ellada"
"Y15-24","EL64",2010,36.9,"Sterea Ellada"
"Y15-24","EL65",2010,29,"Peloponnisos"
"Y15-24","ES",2010,41.5,"Spain"
"Y15-24","ES1",2010,35.9,"Noroeste (ES)"
"Y15-24","ES11",2010,35.4,"Galicia"
"Y15-24","ES12",2010,37.3,"Principado de Asturias"
"Y15-24","ES13",2010,36.1,"Cantabria"
"Y15-24","ES2",2010,31.5,"Noreste (ES)"
"Y15-24","ES21",2010,30.6,"País Vasco"
"Y15-24","ES22",2010,30.4,"Comunidad Foral de Navarra"
"Y15-24","ES23",2010,38.2,"La Rioja"
"Y15-24","ES24",2010,31.9,"Aragón"
"Y15-24","ES3",2010,37.1,"Comunidad de Madrid"
"Y15-24","ES30",2010,37.1,"Comunidad de Madrid"
"Y15-24","ES4",2010,40.2,"Centro (ES)"
"Y15-24","ES41",2010,34,"Castilla y León"
"Y15-24","ES42",2010,42.9,"Castilla-la Mancha"
"Y15-24","ES43",2010,45.8,"Extremadura"
"Y15-24","ES5",2010,40.5,"Este (ES)"
"Y15-24","ES51",2010,39.1,"Cataluña"
"Y15-24","ES52",2010,42.2,"Comunidad Valenciana"
"Y15-24","ES53",2010,42.7,"Illes Balears"
"Y15-24","ES6",2010,48.5,"Sur (ES)"
"Y15-24","ES61",2010,49.9,"Andalucía"
"Y15-24","ES62",2010,39.4,"Región de Murcia"
"Y15-24","ES63",2010,62.1,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2010,52,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2010,52,"Canarias (ES)"
"Y15-24","ES70",2010,52,"Canarias (ES)"
"Y15-24","EU15",2010,20.5,"European Union (15 countries)"
"Y15-24","EU27",2010,21.1,"European Union (27 countries)"
"Y15-24","EU28",2010,21.2,"European Union (28 countries)"
"Y15-24","FI",2010,21.4,"Finland"
"Y15-24","FI1",2010,21.4,"Manner-Suomi"
"Y15-24","FI19",2010,22.8,"Länsi-Suomi"
"Y15-24","FI1B",2010,18.4,"Helsinki-Uusimaa"
"Y15-24","FI1C",2010,21.8,"Etelä-Suomi"
"Y15-24","FI1D",2010,23.9,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2010,NA,"Åland"
"Y15-24","FI20",2010,NA,"Åland"
"Y15-24","FR",2010,23.5,"France"
"Y15-24","FR1",2010,21.2,"Île de France"
"Y15-24","FR10",2010,21.2,"Île de France"
"Y15-24","FR2",2010,23,"Bassin Parisien"
"Y15-24","FR21",2010,24.5,"Champagne-Ardenne"
"Y15-24","FR22",2010,28.2,"Picardie"
"Y15-24","FR23",2010,28.9,"Haute-Normandie"
"Y15-24","FR24",2010,16.2,"Centre (FR)"
"Y15-24","FR25",2010,19.9,"Basse-Normandie"
"Y15-24","FR26",2010,22.6,"Bourgogne"
"Y15-24","FR3",2010,30.1,"Nord - Pas-de-Calais"
"Y15-24","FR30",2010,30.1,"Nord - Pas-de-Calais"
"Y15-24","FR4",2010,21.5,"Est (FR)"
"Y15-24","FR41",2010,24.3,"Lorraine"
"Y15-24","FR42",2010,18.4,"Alsace"
"Y15-24","FR43",2010,20.8,"Franche-Comté"
"Y15-24","FR5",2010,18.7,"Ouest (FR)"
"Y15-24","FR51",2010,18.2,"Pays de la Loire"
"Y15-24","FR52",2010,19,"Bretagne"
"Y15-24","FR53",2010,19.8,"Poitou-Charentes"
"Y15-24","FR6",2010,22.8,"Sud-Ouest (FR)"
"Y15-24","FR61",2010,24.8,"Aquitaine"
"Y15-24","FR62",2010,21.9,"Midi-Pyrénées"
"Y15-24","FR63",2010,18.7,"Limousin"
"Y15-24","FR7",2010,20.2,"Centre-Est (FR)"
"Y15-24","FR71",2010,20.3,"Rhône-Alpes"
"Y15-24","FR72",2010,19.5,"Auvergne"
"Y15-24","FR8",2010,26.6,"Méditerranée"
"Y15-24","FR81",2010,33.2,"Languedoc-Roussillon"
"Y15-24","FR82",2010,23.8,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2010,NA,"Corse"
"Y15-24","FRA",2010,54.2,"Départements d'outre-mer"
"Y15-24","FRA1",2010,55.1,"Guadeloupe"
"Y15-24","FRA2",2010,59,"Martinique"
"Y15-24","FRA3",2010,42.6,"Guyane"
"Y15-24","FRA4",2010,54.7,"La Réunion"
"Y15-24","HR",2010,32.4,"Croatia"
"Y15-24","HR0",2010,32.4,"Hrvatska"
"Y15-24","HR03",2010,27.8,"Jadranska Hrvatska"
"Y15-24","HR04",2010,34.3,"Kontinentalna Hrvatska"
"Y15-24","HU",2010,26.4,"Hungary"
"Y15-24","HU1",2010,21.3,"Közép-Magyarország"
"Y15-24","HU10",2010,21.3,"Közép-Magyarország"
"Y15-24","HU2",2010,24.4,"Dunántúl"
"Y15-24","HU21",2010,21.4,"Közép-Dunántúl"
"Y15-24","HU22",2010,24.4,"Nyugat-Dunántúl"
"Y15-24","HU23",2010,28.3,"Dél-Dunántúl"
"Y15-24","HU3",2010,31,"Alföld és Észak"
"Y15-24","HU31",2010,31.7,"Észak-Magyarország"
"Y15-24","HU32",2010,34.2,"Észak-Alföld"
"Y15-24","HU33",2010,25.7,"Dél-Alföld"
"Y15-24","IE",2010,27.6,"Ireland"
"Y15-24","IE0",2010,27.6,"Éire/Ireland"
"Y15-24","IE01",2010,29.8,"Border, Midland and Western"
"Y15-24","IE02",2010,26.8,"Southern and Eastern"
"Y15-24","IS",2010,16.2,"Iceland"
"Y15-24","IS0",2010,16.2,"Ísland"
"Y15-24","IS00",2010,16.2,"Ísland"
"Y15-24","IT",2010,27.9,"Italy"
"Y15-24","ITC",2010,22,"Nord-Ovest"
"Y15-24","ITC1",2010,26.6,"Piemonte"
"Y15-24","ITC2",2010,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2010,21.3,"Liguria"
"Y15-24","ITC4",2010,20,"Lombardia"
"Y15-24","ITF",2010,37.7,"Sud"
"Y15-24","ITF1",2010,29.5,"Abruzzo"
"Y15-24","ITF2",2010,30.6,"Molise"
"Y15-24","ITF3",2010,41.8,"Campania"
"Y15-24","ITF4",2010,34.6,"Puglia"
"Y15-24","ITF5",2010,41.7,"Basilicata"
"Y15-24","ITF6",2010,38.8,"Calabria"
"Y15-24","ITG",2010,40.9,"Isole"
"Y15-24","ITG1",2010,41.7,"Sicilia"
"Y15-24","ITG2",2010,38.6,"Sardegna"
"Y15-24","ITH",2010,18.8,"Nord-Est"
"Y15-24","ITH1",2010,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2010,15.1,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2010,18.8,"Veneto"
"Y15-24","ITH4",2010,17.6,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2010,22.2,"Emilia-Romagna"
"Y15-24","ITI",2010,25.6,"Centro (IT)"
"Y15-24","ITI1",2010,23,"Toscana"
"Y15-24","ITI2",2010,21.4,"Umbria"
"Y15-24","ITI3",2010,15.2,"Marche"
"Y15-24","ITI4",2010,30.9,"Lazio"
"Y15-24","LT",2010,35.7,"Lithuania"
"Y15-24","LT0",2010,35.7,"Lietuva"
"Y15-24","LT00",2010,35.7,"Lietuva"
"Y15-24","LU",2010,14.2,"Luxembourg"
"Y15-24","LU0",2010,14.2,"Luxembourg"
"Y15-24","LU00",2010,14.2,"Luxembourg"
"Y15-24","LV",2010,36.2,"Latvia"
"Y15-24","LV0",2010,36.2,"Latvija"
"Y15-24","LV00",2010,36.2,"Latvija"
"Y15-24","MK",2010,53.7,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2010,53.7,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2010,53.7,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2010,13.2,"Malta"
"Y15-24","MT0",2010,13.2,"Malta"
"Y15-24","MT00",2010,13.2,"Malta"
"Y15-24","NL",2010,8.7,"Netherlands"
"Y15-24","NL1",2010,9.2,"Noord-Nederland"
"Y15-24","NL11",2010,9.6,"Groningen"
"Y15-24","NL12",2010,9,"Friesland (NL)"
"Y15-24","NL13",2010,9.1,"Drenthe"
"Y15-24","NL2",2010,8.7,"Oost-Nederland"
"Y15-24","NL21",2010,8.5,"Overijssel"
"Y15-24","NL22",2010,8.2,"Gelderland"
"Y15-24","NL23",2010,11.9,"Flevoland"
"Y15-24","NL3",2010,8.8,"West-Nederland"
"Y15-24","NL31",2010,7.1,"Utrecht"
"Y15-24","NL32",2010,8.4,"Noord-Holland"
"Y15-24","NL33",2010,10.2,"Zuid-Holland"
"Y15-24","NL34",2010,NA,"Zeeland"
"Y15-24","NL4",2010,8.1,"Zuid-Nederland"
"Y15-24","NL41",2010,7.5,"Noord-Brabant"
"Y15-24","NL42",2010,9.5,"Limburg (NL)"
"Y15-24","NO",2010,9.3,"Norway"
"Y15-24","NO0",2010,9.3,"Norge"
"Y15-24","NO01",2010,10.1,"Oslo og Akershus"
"Y15-24","NO02",2010,11.1,"Hedmark og Oppland"
"Y15-24","NO03",2010,9.6,"Sør-Østlandet"
"Y15-24","NO04",2010,5.6,"Agder og Rogaland"
"Y15-24","NO05",2010,8.8,"Vestlandet"
"Y15-24","NO06",2010,10.1,"Trøndelag"
"Y15-24","NO07",2010,11.4,"Nord-Norge"
"Y15-24","PL",2010,23.7,"Poland"
"Y15-24","PL1",2010,19.8,"Region Centralny"
"Y15-24","PL11",2010,21.3,"Lódzkie"
"Y15-24","PL12",2010,19.1,"Mazowieckie"
"Y15-24","PL2",2010,22.9,"Region Poludniowy"
"Y15-24","PL21",2010,21.5,"Malopolskie"
"Y15-24","PL22",2010,24,"Slaskie"
"Y15-24","PL3",2010,29.1,"Region Wschodni"
"Y15-24","PL31",2010,26.1,"Lubelskie"
"Y15-24","PL32",2010,35.3,"Podkarpackie"
"Y15-24","PL33",2010,28.2,"Swietokrzyskie"
"Y15-24","PL34",2010,24.5,"Podlaskie"
"Y15-24","PL4",2010,24,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2010,21.8,"Wielkopolskie"
"Y15-24","PL42",2010,30.9,"Zachodniopomorskie"
"Y15-24","PL43",2010,24.3,"Lubuskie"
"Y15-24","PL5",2010,23.2,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2010,23.8,"Dolnoslaskie"
"Y15-24","PL52",2010,21.5,"Opolskie"
"Y15-24","PL6",2010,23.4,"Region Pólnocny"
"Y15-24","PL61",2010,25.4,"Kujawsko-Pomorskie"
"Y15-24","PL62",2010,24,"Warminsko-Mazurskie"
"Y15-24","PL63",2010,21,"Pomorskie"
"Y15-24","PT",2010,22.8,"Portugal"
"Y15-24","PT1",2010,23.1,"Continente"
"Y15-24","PT11",2010,23.2,"Norte"
"Y15-24","PT15",2010,28.9,"Algarve"
"Y15-24","PT16",2010,17.7,"Centro (PT)"
"Y15-24","PT17",2010,25,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2010,29.5,"Alentejo"
"Y15-24","PT2",2010,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2010,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2010,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2010,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2010,22.1,"Romania"
"Y15-24","RO1",2010,25.1,"Macroregiunea unu"
"Y15-24","RO11",2010,18.9,"Nord-Vest"
"Y15-24","RO12",2010,33.2,"Centru"
"Y15-24","RO2",2010,18.2,"Macroregiunea doi"
"Y15-24","RO21",2010,13.5,"Nord-Est"
"Y15-24","RO22",2010,26.1,"Sud-Est"
"Y15-24","RO3",2010,25.9,"Macroregiunea trei"
"Y15-24","RO31",2010,29.2,"Sud - Muntenia"
"Y15-24","RO32",2010,20.1,"Bucuresti - Ilfov"
"Y15-24","RO4",2010,19.2,"Macroregiunea patru"
"Y15-24","RO41",2010,18.6,"Sud-Vest Oltenia"
"Y15-24","RO42",2010,20.1,"Vest"
"Y15-24","SE",2010,24.8,"Sweden"
"Y15-24","SE1",2010,23.5,"Östra Sverige"
"Y15-24","SE11",2010,21,"Stockholm"
"Y15-24","SE12",2010,26.5,"Östra Mellansverige"
"Y15-24","SE2",2010,24.9,"Södra Sverige"
"Y15-24","SE21",2010,21.6,"Småland med öarna"
"Y15-24","SE22",2010,26.7,"Sydsverige"
"Y15-24","SE23",2010,25.1,"Västsverige"
"Y15-24","SE3",2010,27,"Norra Sverige"
"Y15-24","SE31",2010,24.9,"Norra Mellansverige"
"Y15-24","SE32",2010,32.4,"Mellersta Norrland"
"Y15-24","SE33",2010,26.7,"Övre Norrland"
"Y15-24","SI",2010,14.7,"Slovenia"
"Y15-24","SI0",2010,14.7,"Slovenija"
"Y15-24","SI03",2010,15.4,"Vzhodna Slovenija"
"Y15-24","SI04",2010,13.9,"Zahodna Slovenija"
"Y15-24","SK",2010,33.6,"Slovakia"
"Y15-24","SK0",2010,33.6,"Slovensko"
"Y15-24","SK01",2010,15.2,"Bratislavský kraj"
"Y15-24","SK02",2010,30.8,"Západné Slovensko"
"Y15-24","SK03",2010,36.2,"Stredné Slovensko"
"Y15-24","SK04",2010,39.7,"Východné Slovensko"
"Y15-24","TR",2010,19.7,"Turkey"
"Y15-24","TR1",2010,21.9,"Istanbul"
"Y15-24","TR10",2010,21.9,"Istanbul"
"Y15-24","TR2",2010,15.5,"Bati Marmara"
"Y15-24","TR21",2010,18.2,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2010,12.2,"Balikesir, Çanakkale"
"Y15-24","TR3",2010,22,"Ege"
"Y15-24","TR31",2010,26.8,"Izmir"
"Y15-24","TR32",2010,19.9,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2010,16.3,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2010,19.2,"Dogu Marmara"
"Y15-24","TR41",2010,17.5,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2010,20.8,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2010,19.3,"Bati Anadolu"
"Y15-24","TR51",2010,23.2,"Ankara"
"Y15-24","TR52",2010,13.6,"Konya, Karaman"
"Y15-24","TR6",2010,21.7,"Akdeniz"
"Y15-24","TR61",2010,19.9,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2010,24.5,"Adana, Mersin"
"Y15-24","TR63",2010,19.1,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2010,21.2,"Orta Anadolu"
"Y15-24","TR71",2010,17.4,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2010,23.7,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2010,14.9,"Bati Karadeniz"
"Y15-24","TR81",2010,27.9,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2010,14,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2010,10.4,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2010,15.3,"Dogu Karadeniz"
"Y15-24","TR90",2010,15.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2010,13.6,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2010,12.3,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2010,14.7,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2010,24.4,"Ortadogu Anadolu"
"Y15-24","TRB1",2010,22.8,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2010,25.7,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2010,15.4,"Güneydogu Anadolu"
"Y15-24","TRC1",2010,16.9,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2010,13.6,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2010,16.2,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2010,19.9,"United Kingdom"
"Y15-24","UKC",2010,20.9,"North East (UK)"
"Y15-24","UKC1",2010,20.3,"Tees Valley and Durham"
"Y15-24","UKC2",2010,21.4,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2010,20.7,"North West (UK)"
"Y15-24","UKD1",2010,24.7,"Cumbria"
"Y15-24","UKD3",2010,22.1,"Greater Manchester"
"Y15-24","UKD4",2010,15.6,"Lancashire"
"Y15-24","UKD6",2010,15.9,"Cheshire"
"Y15-24","UKD7",2010,24.6,"Merseyside"
"Y15-24","UKE",2010,21.2,"Yorkshire and The Humber"
"Y15-24","UKE1",2010,23.2,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2010,20.3,"North Yorkshire"
"Y15-24","UKE3",2010,20.1,"South Yorkshire"
"Y15-24","UKE4",2010,21.2,"West Yorkshire"
"Y15-24","UKF",2010,18.5,"East Midlands (UK)"
"Y15-24","UKF1",2010,21.3,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2010,18,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2010,11.3,"Lincolnshire"
"Y15-24","UKG",2010,22.7,"West Midlands (UK)"
"Y15-24","UKG1",2010,22,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2010,18.2,"Shropshire and Staffordshire"
"Y15-24","UKG3",2010,25.5,"West Midlands"
"Y15-24","UKH",2010,17.2,"East of England"
"Y15-24","UKH1",2010,18.2,"East Anglia"
"Y15-24","UKH2",2010,17,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2010,16,"Essex"
"Y15-24","UKI",2010,23.9,"London"
"Y15-24","UKI3",2010,20.9,"Inner London - West"
"Y15-24","UKI4",2010,28.9,"Inner London - East"
"Y15-24","UKI5",2010,24.2,"Outer London - East and North East"
"Y15-24","UKI6",2010,18.5,"Outer London - South"
"Y15-24","UKI7",2010,22,"Outer London - West and North West"
"Y15-24","UKJ",2010,16.3,"South East (UK)"
"Y15-24","UKJ1",2010,13.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2010,13.8,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2010,17.3,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2010,21.6,"Kent"
"Y15-24","UKK",2010,15.6,"South West (UK)"
"Y15-24","UKK1",2010,14.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2010,11.6,"Dorset and Somerset"
"Y15-24","UKK3",2010,24.2,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2010,18.5,"Devon"
"Y15-24","UKL",2010,24.6,"Wales"
"Y15-24","UKL1",2010,26.8,"West Wales and The Valleys"
"Y15-24","UKL2",2010,21,"East Wales"
"Y15-24","UKM",2010,19.7,"Scotland"
"Y15-24","UKM2",2010,19.8,"Eastern Scotland"
"Y15-24","UKM3",2010,21.6,"South Western Scotland"
"Y15-24","UKM5",2010,12.4,"North Eastern Scotland"
"Y15-24","UKM6",2010,19.2,"Highlands and Islands"
"Y15-24","UKN",2010,19,"Northern Ireland (UK)"
"Y15-24","UKN0",2010,19,"Northern Ireland (UK)"
"Y20-64","AT",2010,4.6,"Austria"
"Y20-64","AT1",2010,5.8,"Ostösterreich"
"Y20-64","AT11",2010,3.5,"Burgenland (AT)"
"Y20-64","AT12",2010,3.8,"Niederösterreich"
"Y20-64","AT13",2010,8.1,"Wien"
"Y20-64","AT2",2010,4.2,"Südösterreich"
"Y20-64","AT21",2010,4.2,"Kärnten"
"Y20-64","AT22",2010,4.2,"Steiermark"
"Y20-64","AT3",2010,3.4,"Westösterreich"
"Y20-64","AT31",2010,3.7,"Oberösterreich"
"Y20-64","AT32",2010,2.9,"Salzburg"
"Y20-64","AT33",2010,2.8,"Tirol"
"Y20-64","AT34",2010,4.1,"Vorarlberg"
"Y20-64","BE",2010,8,"Belgium"
"Y20-64","BE1",2010,17,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2010,17,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2010,4.9,"Vlaams Gewest"
"Y20-64","BE21",2010,5.8,"Prov. Antwerpen"
"Y20-64","BE22",2010,5,"Prov. Limburg (BE)"
"Y20-64","BE23",2010,5,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2010,4.6,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2010,3.7,"Prov. West-Vlaanderen"
"Y20-64","BE3",2010,11,"Région wallonne"
"Y20-64","BE31",2010,7.8,"Prov. Brabant Wallon"
"Y20-64","BE32",2010,13.3,"Prov. Hainaut"
"Y20-64","BE33",2010,11.2,"Prov. Liège"
"Y20-64","BE34",2010,7.2,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2010,9.5,"Prov. Namur"
"Y20-64","BG",2010,10,"Bulgaria"
"Y20-64","BG3",2010,11.8,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2010,10.9,"Severozapaden"
"Y20-64","BG32",2010,11.4,"Severen tsentralen"
"Y20-64","BG33",2010,14.4,"Severoiztochen"
"Y20-64","BG34",2010,10.2,"Yugoiztochen"
"Y20-64","BG4",2010,8.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2010,6.7,"Yugozapaden"
"Y20-64","BG42",2010,11.1,"Yuzhen tsentralen"
"Y20-64","CH",2010,4.5,"Switzerland"
"Y20-64","CH0",2010,4.5,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2010,6.3,"Région lémanique"
"Y20-64","CH02",2010,4.2,"Espace Mittelland"
"Y20-64","CH03",2010,4.5,"Nordwestschweiz"
"Y20-64","CH04",2010,4.3,"Zürich"
"Y20-64","CH05",2010,3.6,"Ostschweiz"
"Y20-64","CH06",2010,3,"Zentralschweiz"
"Y20-64","CH07",2010,5.9,"Ticino"
"Y20-64","CY",2010,6.2,"Cyprus"
"Y20-64","CY0",2010,6.2,"Kypros"
"Y20-64","CY00",2010,6.2,"Kypros"
"Y20-64","CZ",2010,7.1,"Czech Republic"
"Y20-64","CZ0",2010,7.1,"Ceská republika"
"Y20-64","CZ01",2010,3.6,"Praha"
"Y20-64","CZ02",2010,5.1,"Strední Cechy"
"Y20-64","CZ03",2010,5.4,"Jihozápad"
"Y20-64","CZ04",2010,10.5,"Severozápad"
"Y20-64","CZ05",2010,6.8,"Severovýchod"
"Y20-64","CZ06",2010,7.5,"Jihovýchod"
"Y20-64","CZ07",2010,8.7,"Strední Morava"
"Y20-64","CZ08",2010,10,"Moravskoslezsko"
"Y20-64","DE",2010,7,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2010,4.7,"Baden-Württemberg"
"Y20-64","DE11",2010,5,"Stuttgart"
"Y20-64","DE12",2010,5.2,"Karlsruhe"
"Y20-64","DE13",2010,3.8,"Freiburg"
"Y20-64","DE14",2010,4.5,"Tübingen"
"Y20-64","DE2",2010,4.3,"Bayern"
"Y20-64","DE21",2010,3.6,"Oberbayern"
"Y20-64","DE22",2010,3.9,"Niederbayern"
"Y20-64","DE23",2010,4,"Oberpfalz"
"Y20-64","DE24",2010,5.8,"Oberfranken"
"Y20-64","DE25",2010,5.4,"Mittelfranken"
"Y20-64","DE26",2010,5,"Unterfranken"
"Y20-64","DE27",2010,4.2,"Schwaben"
"Y20-64","DE3",2010,12.9,"Berlin"
"Y20-64","DE30",2010,12.9,"Berlin"
"Y20-64","DE4",2010,9.8,"Brandenburg"
"Y20-64","DE40",2010,9.8,"Brandenburg"
"Y20-64","DE5",2010,8,"Bremen"
"Y20-64","DE50",2010,8,"Bremen"
"Y20-64","DE6",2010,7,"Hamburg"
"Y20-64","DE60",2010,7,"Hamburg"
"Y20-64","DE7",2010,5.7,"Hessen"
"Y20-64","DE71",2010,5.6,"Darmstadt"
"Y20-64","DE72",2010,5.7,"Gießen"
"Y20-64","DE73",2010,5.9,"Kassel"
"Y20-64","DE8",2010,12.4,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2010,12.4,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2010,6.3,"Niedersachsen"
"Y20-64","DE91",2010,7,"Braunschweig"
"Y20-64","DE92",2010,7,"Hannover"
"Y20-64","DE93",2010,5.5,"Lüneburg"
"Y20-64","DE94",2010,5.9,"Weser-Ems"
"Y20-64","DEA",2010,7.3,"Nordrhein-Westfalen"
"Y20-64","DEA1",2010,7.6,"Düsseldorf"
"Y20-64","DEA2",2010,6.9,"Köln"
"Y20-64","DEA3",2010,6.6,"Münster"
"Y20-64","DEA4",2010,6.9,"Detmold"
"Y20-64","DEA5",2010,8.1,"Arnsberg"
"Y20-64","DEB",2010,5.3,"Rheinland-Pfalz"
"Y20-64","DEB1",2010,5.2,"Koblenz"
"Y20-64","DEB2",2010,4,"Trier"
"Y20-64","DEB3",2010,5.8,"Rheinhessen-Pfalz"
"Y20-64","DEC",2010,6.6,"Saarland"
"Y20-64","DEC0",2010,6.6,"Saarland"
"Y20-64","DED",2010,11.3,"Sachsen"
"Y20-64","DED2",2010,10.4,"Dresden"
"Y20-64","DED4",2010,11.7,"Chemnitz"
"Y20-64","DED5",2010,12.3,"Leipzig"
"Y20-64","DEE",2010,11.4,"Sachsen-Anhalt"
"Y20-64","DEE0",2010,11.4,"Sachsen-Anhalt"
"Y20-64","DEF",2010,6.5,"Schleswig-Holstein"
"Y20-64","DEF0",2010,6.5,"Schleswig-Holstein"
"Y20-64","DEG",2010,8.6,"Thüringen"
"Y20-64","DEG0",2010,8.6,"Thüringen"
"Y20-64","DK",2010,6.9,"Denmark"
"Y20-64","DK0",2010,6.9,"Danmark"
"Y20-64","DK01",2010,7.3,"Hovedstaden"
"Y20-64","DK02",2010,6,"Sjælland"
"Y20-64","DK03",2010,7,"Syddanmark"
"Y20-64","DK04",2010,6.7,"Midtjylland"
"Y20-64","DK05",2010,7.2,"Nordjylland"
"Y20-64","EA17",2010,9.8,"Euro area (17 countries)"
"Y20-64","EA18",2010,9.8,"Euro area (18 countries)"
"Y20-64","EA19",2010,9.9,"Euro area (19 countries)"
"Y20-64","EE",2010,16.7,"Estonia"
"Y20-64","EE0",2010,16.7,"Eesti"
"Y20-64","EE00",2010,16.7,"Eesti"
"Y20-64","EL",2010,12.7,"Greece"
"Y20-64","EL3",2010,12.6,"Attiki"
"Y20-64","EL30",2010,12.6,"Attiki"
"Y20-64","EL4",2010,12.2,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2010,9.1,"Voreio Aigaio"
"Y20-64","EL42",2010,14.2,"Notio Aigaio"
"Y20-64","EL43",2010,12,"Kriti"
"Y20-64","EL5",2010,13.8,"Voreia Ellada"
"Y20-64","EL51",2010,14.2,"Anatoliki Makedonia, Thraki"
"Y20-64","EL52",2010,13.6,"Kentriki Makedonia"
"Y20-64","EL53",2010,15.5,"Dytiki Makedonia"
"Y20-64","EL54",2010,12.7,"Ipeiros"
"Y20-64","EL6",2010,11.8,"Kentriki Ellada"
"Y20-64","EL61",2010,12.2,"Thessalia"
"Y20-64","EL62",2010,14.5,"Ionia Nisia"
"Y20-64","EL63",2010,11.8,"Dytiki Ellada"
"Y20-64","EL64",2010,12.2,"Sterea Ellada"
"Y20-64","EL65",2010,9.7,"Peloponnisos"
"Y20-64","ES",2010,19.3,"Spain"
"Y20-64","ES1",2010,14.9,"Noroeste (ES)"
"Y20-64","ES11",2010,15,"Galicia"
"Y20-64","ES12",2010,15.6,"Principado de Asturias"
"Y20-64","ES13",2010,13.4,"Cantabria"
"Y20-64","ES2",2010,12.1,"Noreste (ES)"
"Y20-64","ES21",2010,10.5,"País Vasco"
"Y20-64","ES22",2010,11.5,"Comunidad Foral de Navarra"
"Y20-64","ES23",2010,13.4,"La Rioja"
"Y20-64","ES24",2010,14.6,"Aragón"
"Y20-64","ES3",2010,15.4,"Comunidad de Madrid"
"Y20-64","ES30",2010,15.4,"Comunidad de Madrid"
"Y20-64","ES4",2010,18.6,"Centro (ES)"
"Y20-64","ES41",2010,15.4,"Castilla y León"
"Y20-64","ES42",2010,20.5,"Castilla-la Mancha"
"Y20-64","ES43",2010,22.3,"Extremadura"
"Y20-64","ES5",2010,19,"Este (ES)"
"Y20-64","ES51",2010,16.9,"Cataluña"
"Y20-64","ES52",2010,22.1,"Comunidad Valenciana"
"Y20-64","ES53",2010,19.2,"Illes Balears"
"Y20-64","ES6",2010,26.2,"Sur (ES)"
"Y20-64","ES61",2010,27,"Andalucía"
"Y20-64","ES62",2010,22.3,"Región de Murcia"
"Y20-64","ES63",2010,23.1,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2010,21.5,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2010,28.2,"Canarias (ES)"
"Y20-64","ES70",2010,28.2,"Canarias (ES)"
"Y20-64","EU15",2010,9.1,"European Union (15 countries)"
"Y20-64","EU27",2010,9.3,"European Union (27 countries)"
"Y20-64","EU28",2010,9.3,"European Union (28 countries)"
"Y20-64","FI",2010,7.6,"Finland"
"Y20-64","FI1",2010,7.7,"Manner-Suomi"
"Y20-64","FI19",2010,8.2,"Länsi-Suomi"
"Y20-64","FI1B",2010,5.5,"Helsinki-Uusimaa"
"Y20-64","FI1C",2010,8.4,"Etelä-Suomi"
"Y20-64","FI1D",2010,9.4,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2010,NA,"Åland"
"Y20-64","FI20",2010,NA,"Åland"
"Y20-64","FR",2010,8.9,"France"
"Y20-64","FR1",2010,8.4,"Île de France"
"Y20-64","FR10",2010,8.4,"Île de France"
"Y20-64","FR2",2010,8.4,"Bassin Parisien"
"Y20-64","FR21",2010,8.5,"Champagne-Ardenne"
"Y20-64","FR22",2010,10.8,"Picardie"
"Y20-64","FR23",2010,8.9,"Haute-Normandie"
"Y20-64","FR24",2010,6.6,"Centre (FR)"
"Y20-64","FR25",2010,8,"Basse-Normandie"
"Y20-64","FR26",2010,8.4,"Bourgogne"
"Y20-64","FR3",2010,11.9,"Nord - Pas-de-Calais"
"Y20-64","FR30",2010,11.9,"Nord - Pas-de-Calais"
"Y20-64","FR4",2010,8.3,"Est (FR)"
"Y20-64","FR41",2010,8.9,"Lorraine"
"Y20-64","FR42",2010,7.6,"Alsace"
"Y20-64","FR43",2010,8,"Franche-Comté"
"Y20-64","FR5",2010,7.4,"Ouest (FR)"
"Y20-64","FR51",2010,8.2,"Pays de la Loire"
"Y20-64","FR52",2010,6.5,"Bretagne"
"Y20-64","FR53",2010,7.3,"Poitou-Charentes"
"Y20-64","FR6",2010,7.4,"Sud-Ouest (FR)"
"Y20-64","FR61",2010,7.5,"Aquitaine"
"Y20-64","FR62",2010,7.4,"Midi-Pyrénées"
"Y20-64","FR63",2010,6.9,"Limousin"
"Y20-64","FR7",2010,7.5,"Centre-Est (FR)"
"Y20-64","FR71",2010,7.7,"Rhône-Alpes"
"Y20-64","FR72",2010,6.9,"Auvergne"
"Y20-64","FR8",2010,10.3,"Méditerranée"
"Y20-64","FR81",2010,13,"Languedoc-Roussillon"
"Y20-64","FR82",2010,9.2,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2010,5.8,"Corse"
"Y20-64","FRA",2010,24.5,"Départements d'outre-mer"
"Y20-64","FRA1",2010,23.5,"Guadeloupe"
"Y20-64","FRA2",2010,20.5,"Martinique"
"Y20-64","FRA3",2010,20.5,"Guyane"
"Y20-64","FRA4",2010,27.9,"La Réunion"
"Y20-64","HR",2010,11.1,"Croatia"
"Y20-64","HR0",2010,11.1,"Hrvatska"
"Y20-64","HR03",2010,10.8,"Jadranska Hrvatska"
"Y20-64","HR04",2010,11.3,"Kontinentalna Hrvatska"
"Y20-64","HU",2010,11.1,"Hungary"
"Y20-64","HU1",2010,8.9,"Közép-Magyarország"
"Y20-64","HU10",2010,8.9,"Közép-Magyarország"
"Y20-64","HU2",2010,10.4,"Dunántúl"
"Y20-64","HU21",2010,9.9,"Közép-Dunántúl"
"Y20-64","HU22",2010,9.2,"Nyugat-Dunántúl"
"Y20-64","HU23",2010,12.3,"Dél-Dunántúl"
"Y20-64","HU3",2010,13.4,"Alföld és Észak"
"Y20-64","HU31",2010,16,"Észak-Magyarország"
"Y20-64","HU32",2010,14.2,"Észak-Alföld"
"Y20-64","HU33",2010,10.3,"Dél-Alföld"
"Y20-64","IE",2010,13.6,"Ireland"
"Y20-64","IE0",2010,13.6,"Éire/Ireland"
"Y20-64","IE01",2010,14.2,"Border, Midland and Western"
"Y20-64","IE02",2010,13.4,"Southern and Eastern"
"Y20-64","IS",2010,6.8,"Iceland"
"Y20-64","IS0",2010,6.8,"Ísland"
"Y20-64","IS00",2010,6.8,"Ísland"
"Y20-64","IT",2010,8.1,"Italy"
"Y20-64","ITC",2010,5.9,"Nord-Ovest"
"Y20-64","ITC1",2010,7.2,"Piemonte"
"Y20-64","ITC2",2010,4.4,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2010,6.4,"Liguria"
"Y20-64","ITC4",2010,5.3,"Lombardia"
"Y20-64","ITF",2010,12.4,"Sud"
"Y20-64","ITF1",2010,8.5,"Abruzzo"
"Y20-64","ITF2",2010,8.2,"Molise"
"Y20-64","ITF3",2010,13.7,"Campania"
"Y20-64","ITF4",2010,13,"Puglia"
"Y20-64","ITF5",2010,12.6,"Basilicata"
"Y20-64","ITF6",2010,11.5,"Calabria"
"Y20-64","ITG",2010,14,"Isole"
"Y20-64","ITG1",2010,14.1,"Sicilia"
"Y20-64","ITG2",2010,13.8,"Sardegna"
"Y20-64","ITH",2010,5.2,"Nord-Est"
"Y20-64","ITH1",2010,2.6,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2010,4,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2010,5.3,"Veneto"
"Y20-64","ITH4",2010,5.5,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2010,5.3,"Emilia-Romagna"
"Y20-64","ITI",2010,7.3,"Centro (IT)"
"Y20-64","ITI1",2010,5.9,"Toscana"
"Y20-64","ITI2",2010,6.3,"Umbria"
"Y20-64","ITI3",2010,5.6,"Marche"
"Y20-64","ITI4",2010,8.9,"Lazio"
"Y20-64","LT",2010,17.8,"Lithuania"
"Y20-64","LT0",2010,17.8,"Lietuva"
"Y20-64","LT00",2010,17.8,"Lietuva"
"Y20-64","LU",2010,4.2,"Luxembourg"
"Y20-64","LU0",2010,4.2,"Luxembourg"
"Y20-64","LU00",2010,4.2,"Luxembourg"
"Y20-64","LV",2010,19.3,"Latvia"
"Y20-64","LV0",2010,19.3,"Latvija"
"Y20-64","LV00",2010,19.3,"Latvija"
"Y20-64","MK",2010,31.6,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2010,31.6,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2010,31.6,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2010,6,"Malta"
"Y20-64","MT0",2010,6,"Malta"
"Y20-64","MT00",2010,6,"Malta"
"Y20-64","NL",2010,4,"Netherlands"
"Y20-64","NL1",2010,4.4,"Noord-Nederland"
"Y20-64","NL11",2010,4.7,"Groningen"
"Y20-64","NL12",2010,4.3,"Friesland (NL)"
"Y20-64","NL13",2010,4.1,"Drenthe"
"Y20-64","NL2",2010,3.7,"Oost-Nederland"
"Y20-64","NL21",2010,3.9,"Overijssel"
"Y20-64","NL22",2010,3.6,"Gelderland"
"Y20-64","NL23",2010,4.2,"Flevoland"
"Y20-64","NL3",2010,4,"West-Nederland"
"Y20-64","NL31",2010,3.3,"Utrecht"
"Y20-64","NL32",2010,3.8,"Noord-Holland"
"Y20-64","NL33",2010,4.5,"Zuid-Holland"
"Y20-64","NL34",2010,2.5,"Zeeland"
"Y20-64","NL4",2010,4.1,"Zuid-Nederland"
"Y20-64","NL41",2010,3.9,"Noord-Brabant"
"Y20-64","NL42",2010,4.8,"Limburg (NL)"
"Y20-64","NO",2010,3.1,"Norway"
"Y20-64","NO0",2010,3.1,"Norge"
"Y20-64","NO01",2010,3.5,"Oslo og Akershus"
"Y20-64","NO02",2010,2.9,"Hedmark og Oppland"
"Y20-64","NO03",2010,3.3,"Sør-Østlandet"
"Y20-64","NO04",2010,2.3,"Agder og Rogaland"
"Y20-64","NO05",2010,3.1,"Vestlandet"
"Y20-64","NO06",2010,3.2,"Trøndelag"
"Y20-64","NO07",2010,3.1,"Nord-Norge"
"Y20-64","PL",2010,9.5,"Poland"
"Y20-64","PL1",2010,8,"Region Centralny"
"Y20-64","PL11",2010,9.1,"Lódzkie"
"Y20-64","PL12",2010,7.4,"Mazowieckie"
"Y20-64","PL2",2010,9,"Region Poludniowy"
"Y20-64","PL21",2010,9,"Malopolskie"
"Y20-64","PL22",2010,9.1,"Slaskie"
"Y20-64","PL3",2010,10.9,"Region Wschodni"
"Y20-64","PL31",2010,10,"Lubelskie"
"Y20-64","PL32",2010,11.6,"Podkarpackie"
"Y20-64","PL33",2010,12,"Swietokrzyskie"
"Y20-64","PL34",2010,10,"Podlaskie"
"Y20-64","PL4",2010,9.8,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2010,8.6,"Wielkopolskie"
"Y20-64","PL42",2010,12.2,"Zachodniopomorskie"
"Y20-64","PL43",2010,10.3,"Lubuskie"
"Y20-64","PL5",2010,10.7,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2010,11.1,"Dolnoslaskie"
"Y20-64","PL52",2010,9.5,"Opolskie"
"Y20-64","PL6",2010,9.7,"Region Pólnocny"
"Y20-64","PL61",2010,10.4,"Kujawsko-Pomorskie"
"Y20-64","PL62",2010,9.5,"Warminsko-Mazurskie"
"Y20-64","PL63",2010,9.1,"Pomorskie"
"Y20-64","PT",2010,11.1,"Portugal"
"Y20-64","PT1",2010,11.3,"Continente"
"Y20-64","PT11",2010,12.9,"Norte"
"Y20-64","PT15",2010,13.4,"Algarve"
"Y20-64","PT16",2010,8.3,"Centro (PT)"
"Y20-64","PT17",2010,11.3,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2010,11.4,"Alentejo"
"Y20-64","PT2",2010,6.5,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2010,6.5,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2010,7.5,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2010,7.5,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2010,7,"Romania"
"Y20-64","RO1",2010,8.1,"Macroregiunea unu"
"Y20-64","RO11",2010,6.6,"Nord-Vest"
"Y20-64","RO12",2010,10,"Centru"
"Y20-64","RO2",2010,6.7,"Macroregiunea doi"
"Y20-64","RO21",2010,5.7,"Nord-Est"
"Y20-64","RO22",2010,8.1,"Sud-Est"
"Y20-64","RO3",2010,6.3,"Macroregiunea trei"
"Y20-64","RO31",2010,7.7,"Sud - Muntenia"
"Y20-64","RO32",2010,4.5,"Bucuresti - Ilfov"
"Y20-64","RO4",2010,6.9,"Macroregiunea patru"
"Y20-64","RO41",2010,7.9,"Sud-Vest Oltenia"
"Y20-64","RO42",2010,5.9,"Vest"
"Y20-64","SE",2010,7.6,"Sweden"
"Y20-64","SE1",2010,7.3,"Östra Sverige"
"Y20-64","SE11",2010,6.3,"Stockholm"
"Y20-64","SE12",2010,8.7,"Östra Mellansverige"
"Y20-64","SE2",2010,7.6,"Södra Sverige"
"Y20-64","SE21",2010,7.1,"Småland med öarna"
"Y20-64","SE22",2010,7.8,"Sydsverige"
"Y20-64","SE23",2010,7.6,"Västsverige"
"Y20-64","SE3",2010,8.4,"Norra Sverige"
"Y20-64","SE31",2010,8.2,"Norra Mellansverige"
"Y20-64","SE32",2010,9.1,"Mellersta Norrland"
"Y20-64","SE33",2010,8.4,"Övre Norrland"
"Y20-64","SI",2010,7.3,"Slovenia"
"Y20-64","SI0",2010,7.3,"Slovenija"
"Y20-64","SI03",2010,7.9,"Vzhodna Slovenija"
"Y20-64","SI04",2010,6.6,"Zahodna Slovenija"
"Y20-64","SK",2010,14,"Slovakia"
"Y20-64","SK0",2010,14,"Slovensko"
"Y20-64","SK01",2010,6.1,"Bratislavský kraj"
"Y20-64","SK02",2010,12.3,"Západné Slovensko"
"Y20-64","SK03",2010,16,"Stredné Slovensko"
"Y20-64","SK04",2010,18,"Východné Slovensko"
"Y20-64","TR",2010,10.5,"Turkey"
"Y20-64","TR1",2010,13.2,"Istanbul"
"Y20-64","TR10",2010,13.2,"Istanbul"
"Y20-64","TR2",2010,7,"Bati Marmara"
"Y20-64","TR21",2010,7.9,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2010,6.2,"Balikesir, Çanakkale"
"Y20-64","TR3",2010,10.7,"Ege"
"Y20-64","TR31",2010,13.8,"Izmir"
"Y20-64","TR32",2010,10.2,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2010,6.7,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2010,9.8,"Dogu Marmara"
"Y20-64","TR41",2010,9,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2010,10.8,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2010,9.2,"Bati Anadolu"
"Y20-64","TR51",2010,10.2,"Ankara"
"Y20-64","TR52",2010,7,"Konya, Karaman"
"Y20-64","TR6",2010,12.1,"Akdeniz"
"Y20-64","TR61",2010,9.5,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2010,14.6,"Adana, Mersin"
"Y20-64","TR63",2010,11.6,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2010,10.9,"Orta Anadolu"
"Y20-64","TR71",2010,9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2010,12.2,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2010,7.6,"Bati Karadeniz"
"Y20-64","TR81",2010,10.3,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2010,7.9,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2010,6.3,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2010,5,"Dogu Karadeniz"
"Y20-64","TR90",2010,5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2010,6.9,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2010,5.7,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2010,8.3,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2010,12.4,"Ortadogu Anadolu"
"Y20-64","TRB1",2010,10.4,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2010,14.7,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2010,10.7,"Güneydogu Anadolu"
"Y20-64","TRC1",2010,11,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2010,11.1,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2010,9.7,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2010,6.8,"United Kingdom"
"Y20-64","UKC",2010,8.3,"North East (UK)"
"Y20-64","UKC1",2010,7.8,"Tees Valley and Durham"
"Y20-64","UKC2",2010,8.8,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2010,6.9,"North West (UK)"
"Y20-64","UKD1",2010,5.5,"Cumbria"
"Y20-64","UKD3",2010,7.5,"Greater Manchester"
"Y20-64","UKD4",2010,5.1,"Lancashire"
"Y20-64","UKD6",2010,4.9,"Cheshire"
"Y20-64","UKD7",2010,9.3,"Merseyside"
"Y20-64","UKE",2010,8,"Yorkshire and The Humber"
"Y20-64","UKE1",2010,7.7,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2010,6.4,"North Yorkshire"
"Y20-64","UKE3",2010,8.4,"South Yorkshire"
"Y20-64","UKE4",2010,8.4,"West Yorkshire"
"Y20-64","UKF",2010,6.7,"East Midlands (UK)"
"Y20-64","UKF1",2010,7.6,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2010,6.4,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2010,4.6,"Lincolnshire"
"Y20-64","UKG",2010,7.8,"West Midlands (UK)"
"Y20-64","UKG1",2010,4.9,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2010,6.7,"Shropshire and Staffordshire"
"Y20-64","UKG3",2010,9.9,"West Midlands"
"Y20-64","UKH",2010,5.7,"East of England"
"Y20-64","UKH1",2010,5.5,"East Anglia"
"Y20-64","UKH2",2010,5.2,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2010,6.6,"Essex"
"Y20-64","UKI",2010,8.2,"London"
"Y20-64","UKI3",2010,7.4,"Inner London - West"
"Y20-64","UKI4",2010,9.9,"Inner London - East"
"Y20-64","UKI5",2010,8.9,"Outer London - East and North East"
"Y20-64","UKI6",2010,6.1,"Outer London - South"
"Y20-64","UKI7",2010,7.7,"Outer London - West and North West"
"Y20-64","UKJ",2010,5.2,"South East (UK)"
"Y20-64","UKJ1",2010,5.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2010,4.5,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2010,5.3,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2010,6.4,"Kent"
"Y20-64","UKK",2010,5.1,"South West (UK)"
"Y20-64","UKK1",2010,4.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2010,4.9,"Dorset and Somerset"
"Y20-64","UKK3",2010,6.6,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2010,5.6,"Devon"
"Y20-64","UKL",2010,7.4,"Wales"
"Y20-64","UKL1",2010,7.9,"West Wales and The Valleys"
"Y20-64","UKL2",2010,6.7,"East Wales"
"Y20-64","UKM",2010,7.2,"Scotland"
"Y20-64","UKM2",2010,6.6,"Eastern Scotland"
"Y20-64","UKM3",2010,9,"South Western Scotland"
"Y20-64","UKM5",2010,2.7,"North Eastern Scotland"
"Y20-64","UKM6",2010,6.2,"Highlands and Islands"
"Y20-64","UKN",2010,6.5,"Northern Ireland (UK)"
"Y20-64","UKN0",2010,6.5,"Northern Ireland (UK)"
"Y_GE15","AT",2010,4.8,"Austria"
"Y_GE15","AT1",2010,6,"Ostösterreich"
"Y_GE15","AT11",2010,4,"Burgenland (AT)"
"Y_GE15","AT12",2010,3.9,"Niederösterreich"
"Y_GE15","AT13",2010,8.3,"Wien"
"Y_GE15","AT2",2010,4.4,"Südösterreich"
"Y_GE15","AT21",2010,4.3,"Kärnten"
"Y_GE15","AT22",2010,4.5,"Steiermark"
"Y_GE15","AT3",2010,3.7,"Westösterreich"
"Y_GE15","AT31",2010,3.9,"Oberösterreich"
"Y_GE15","AT32",2010,3.2,"Salzburg"
"Y_GE15","AT33",2010,3.2,"Tirol"
"Y_GE15","AT34",2010,4.6,"Vorarlberg"
"Y_GE15","BE",2010,8.3,"Belgium"
"Y_GE15","BE1",2010,17.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2010,17.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2010,5.1,"Vlaams Gewest"
"Y_GE15","BE21",2010,6,"Prov. Antwerpen"
"Y_GE15","BE22",2010,5.3,"Prov. Limburg (BE)"
"Y_GE15","BE23",2010,5.2,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2010,4.8,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2010,3.8,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2010,11.4,"Région wallonne"
"Y_GE15","BE31",2010,8.3,"Prov. Brabant Wallon"
"Y_GE15","BE32",2010,13.9,"Prov. Hainaut"
"Y_GE15","BE33",2010,11.5,"Prov. Liège"
"Y_GE15","BE34",2010,7.5,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2010,9.6,"Prov. Namur"
"Y_GE15","BG",2010,10.3,"Bulgaria"
"Y_GE15","BG3",2010,12,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2010,11.2,"Severozapaden"
"Y_GE15","BG32",2010,11.6,"Severen tsentralen"
"Y_GE15","BG33",2010,14.6,"Severoiztochen"
"Y_GE15","BG34",2010,10.5,"Yugoiztochen"
"Y_GE15","BG4",2010,8.7,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2010,6.9,"Yugozapaden"
"Y_GE15","BG42",2010,11.5,"Yuzhen tsentralen"
"Y_GE15","CH",2010,4.5,"Switzerland"
"Y_GE15","CH0",2010,4.5,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2010,6.7,"Région lémanique"
"Y_GE15","CH02",2010,4.2,"Espace Mittelland"
"Y_GE15","CH03",2010,4.5,"Nordwestschweiz"
"Y_GE15","CH04",2010,4.2,"Zürich"
"Y_GE15","CH05",2010,3.5,"Ostschweiz"
"Y_GE15","CH06",2010,3,"Zentralschweiz"
"Y_GE15","CH07",2010,6,"Ticino"
"Y_GE15","CY",2010,6.3,"Cyprus"
"Y_GE15","CY0",2010,6.3,"Kypros"
"Y_GE15","CY00",2010,6.3,"Kypros"
"Y_GE15","CZ",2010,7.3,"Czech Republic"
"Y_GE15","CZ0",2010,7.3,"Ceská republika"
"Y_GE15","CZ01",2010,3.7,"Praha"
"Y_GE15","CZ02",2010,5.2,"Strední Cechy"
"Y_GE15","CZ03",2010,5.6,"Jihozápad"
"Y_GE15","CZ04",2010,11.1,"Severozápad"
"Y_GE15","CZ05",2010,7,"Severovýchod"
"Y_GE15","CZ06",2010,7.5,"Jihovýchod"
"Y_GE15","CZ07",2010,8.8,"Strední Morava"
"Y_GE15","CZ08",2010,10.2,"Moravskoslezsko"
"Y_GE15","DE",2010,7,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2010,4.7,"Baden-Württemberg"
"Y_GE15","DE11",2010,5,"Stuttgart"
"Y_GE15","DE12",2010,5.2,"Karlsruhe"
"Y_GE15","DE13",2010,3.9,"Freiburg"
"Y_GE15","DE14",2010,4.5,"Tübingen"
"Y_GE15","DE2",2010,4.3,"Bayern"
"Y_GE15","DE21",2010,3.6,"Oberbayern"
"Y_GE15","DE22",2010,3.9,"Niederbayern"
"Y_GE15","DE23",2010,4,"Oberpfalz"
"Y_GE15","DE24",2010,5.9,"Oberfranken"
"Y_GE15","DE25",2010,5.5,"Mittelfranken"
"Y_GE15","DE26",2010,5.1,"Unterfranken"
"Y_GE15","DE27",2010,4.2,"Schwaben"
"Y_GE15","DE3",2010,12.8,"Berlin"
"Y_GE15","DE30",2010,12.8,"Berlin"
"Y_GE15","DE4",2010,9.8,"Brandenburg"
"Y_GE15","DE40",2010,9.8,"Brandenburg"
"Y_GE15","DE5",2010,7.9,"Bremen"
"Y_GE15","DE50",2010,7.9,"Bremen"
"Y_GE15","DE6",2010,7,"Hamburg"
"Y_GE15","DE60",2010,7,"Hamburg"
"Y_GE15","DE7",2010,5.9,"Hessen"
"Y_GE15","DE71",2010,5.8,"Darmstadt"
"Y_GE15","DE72",2010,6,"Gießen"
"Y_GE15","DE73",2010,6,"Kassel"
"Y_GE15","DE8",2010,12.3,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2010,12.3,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2010,6.4,"Niedersachsen"
"Y_GE15","DE91",2010,7.1,"Braunschweig"
"Y_GE15","DE92",2010,7,"Hannover"
"Y_GE15","DE93",2010,5.7,"Lüneburg"
"Y_GE15","DE94",2010,5.9,"Weser-Ems"
"Y_GE15","DEA",2010,7.4,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2010,7.6,"Düsseldorf"
"Y_GE15","DEA2",2010,7,"Köln"
"Y_GE15","DEA3",2010,6.6,"Münster"
"Y_GE15","DEA4",2010,7,"Detmold"
"Y_GE15","DEA5",2010,8.2,"Arnsberg"
"Y_GE15","DEB",2010,5.5,"Rheinland-Pfalz"
"Y_GE15","DEB1",2010,5.1,"Koblenz"
"Y_GE15","DEB2",2010,4.1,"Trier"
"Y_GE15","DEB3",2010,6,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2010,6.9,"Saarland"
"Y_GE15","DEC0",2010,6.9,"Saarland"
"Y_GE15","DED",2010,11.2,"Sachsen"
"Y_GE15","DED2",2010,10.3,"Dresden"
"Y_GE15","DED4",2010,11.5,"Chemnitz"
"Y_GE15","DED5",2010,12.1,"Leipzig"
"Y_GE15","DEE",2010,11.4,"Sachsen-Anhalt"
"Y_GE15","DEE0",2010,11.4,"Sachsen-Anhalt"
"Y_GE15","DEF",2010,6.6,"Schleswig-Holstein"
"Y_GE15","DEF0",2010,6.6,"Schleswig-Holstein"
"Y_GE15","DEG",2010,8.6,"Thüringen"
"Y_GE15","DEG0",2010,8.6,"Thüringen"
"Y_GE15","DK",2010,7.5,"Denmark"
"Y_GE15","DK0",2010,7.5,"Danmark"
"Y_GE15","DK01",2010,7.9,"Hovedstaden"
"Y_GE15","DK02",2010,6.8,"Sjælland"
"Y_GE15","DK03",2010,7.6,"Syddanmark"
"Y_GE15","DK04",2010,7.2,"Midtjylland"
"Y_GE15","DK05",2010,7.4,"Nordjylland"
"Y_GE15","EA17",2010,10,"Euro area (17 countries)"
"Y_GE15","EA18",2010,10.1,"Euro area (18 countries)"
"Y_GE15","EA19",2010,10.1,"Euro area (19 countries)"
"Y_GE15","EE",2010,16.7,"Estonia"
"Y_GE15","EE0",2010,16.7,"Eesti"
"Y_GE15","EE00",2010,16.7,"Eesti"
"Y_GE15","EL",2010,12.7,"Greece"
"Y_GE15","EL3",2010,12.6,"Attiki"
"Y_GE15","EL30",2010,12.6,"Attiki"
"Y_GE15","EL4",2010,12.3,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2010,9.4,"Voreio Aigaio"
"Y_GE15","EL42",2010,14.6,"Notio Aigaio"
"Y_GE15","EL43",2010,12,"Kriti"
"Y_GE15","EL5",2010,13.9,"Voreia Ellada"
"Y_GE15","EL51",2010,14.5,"Anatoliki Makedonia, Thraki"
"Y_GE15","EL52",2010,13.7,"Kentriki Makedonia"
"Y_GE15","EL53",2010,15.4,"Dytiki Makedonia"
"Y_GE15","EL54",2010,12.6,"Ipeiros"
"Y_GE15","EL6",2010,11.8,"Kentriki Ellada"
"Y_GE15","EL61",2010,12.1,"Thessalia"
"Y_GE15","EL62",2010,14.6,"Ionia Nisia"
"Y_GE15","EL63",2010,11.9,"Dytiki Ellada"
"Y_GE15","EL64",2010,12.5,"Sterea Ellada"
"Y_GE15","EL65",2010,9.6,"Peloponnisos"
"Y_GE15","ES",2010,19.9,"Spain"
"Y_GE15","ES1",2010,15.2,"Noroeste (ES)"
"Y_GE15","ES11",2010,15.3,"Galicia"
"Y_GE15","ES12",2010,15.9,"Principado de Asturias"
"Y_GE15","ES13",2010,13.7,"Cantabria"
"Y_GE15","ES2",2010,12.4,"Noreste (ES)"
"Y_GE15","ES21",2010,10.7,"País Vasco"
"Y_GE15","ES22",2010,11.9,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2010,14.1,"La Rioja"
"Y_GE15","ES24",2010,15,"Aragón"
"Y_GE15","ES3",2010,15.8,"Comunidad de Madrid"
"Y_GE15","ES30",2010,15.8,"Comunidad de Madrid"
"Y_GE15","ES4",2010,19.1,"Centro (ES)"
"Y_GE15","ES41",2010,15.8,"Castilla y León"
"Y_GE15","ES42",2010,21.2,"Castilla-la Mancha"
"Y_GE15","ES43",2010,23,"Extremadura"
"Y_GE15","ES5",2010,19.7,"Este (ES)"
"Y_GE15","ES51",2010,17.7,"Cataluña"
"Y_GE15","ES52",2010,22.9,"Comunidad Valenciana"
"Y_GE15","ES53",2010,20.1,"Illes Balears"
"Y_GE15","ES6",2010,27,"Sur (ES)"
"Y_GE15","ES61",2010,27.8,"Andalucía"
"Y_GE15","ES62",2010,22.9,"Región de Murcia"
"Y_GE15","ES63",2010,23.9,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2010,22.8,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2010,28.6,"Canarias (ES)"
"Y_GE15","ES70",2010,28.6,"Canarias (ES)"
"Y_GE15","EU15",2010,9.5,"European Union (15 countries)"
"Y_GE15","EU27",2010,9.6,"European Union (27 countries)"
"Y_GE15","EU28",2010,9.6,"European Union (28 countries)"
"Y_GE15","FI",2010,8.4,"Finland"
"Y_GE15","FI1",2010,8.4,"Manner-Suomi"
"Y_GE15","FI19",2010,9,"Länsi-Suomi"
"Y_GE15","FI1B",2010,6.4,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2010,9.1,"Etelä-Suomi"
"Y_GE15","FI1D",2010,10.1,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2010,NA,"Åland"
"Y_GE15","FI20",2010,NA,"Åland"
"Y_GE15","FR",2010,9.3,"France"
"Y_GE15","FR1",2010,8.5,"Île de France"
"Y_GE15","FR10",2010,8.5,"Île de France"
"Y_GE15","FR2",2010,9,"Bassin Parisien"
"Y_GE15","FR21",2010,9.2,"Champagne-Ardenne"
"Y_GE15","FR22",2010,11.4,"Picardie"
"Y_GE15","FR23",2010,9.7,"Haute-Normandie"
"Y_GE15","FR24",2010,7,"Centre (FR)"
"Y_GE15","FR25",2010,8.2,"Basse-Normandie"
"Y_GE15","FR26",2010,8.9,"Bourgogne"
"Y_GE15","FR3",2010,12.5,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2010,12.5,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2010,8.7,"Est (FR)"
"Y_GE15","FR41",2010,9.4,"Lorraine"
"Y_GE15","FR42",2010,8.1,"Alsace"
"Y_GE15","FR43",2010,8.2,"Franche-Comté"
"Y_GE15","FR5",2010,7.7,"Ouest (FR)"
"Y_GE15","FR51",2010,8.5,"Pays de la Loire"
"Y_GE15","FR52",2010,6.8,"Bretagne"
"Y_GE15","FR53",2010,7.7,"Poitou-Charentes"
"Y_GE15","FR6",2010,7.9,"Sud-Ouest (FR)"
"Y_GE15","FR61",2010,8.1,"Aquitaine"
"Y_GE15","FR62",2010,7.8,"Midi-Pyrénées"
"Y_GE15","FR63",2010,7,"Limousin"
"Y_GE15","FR7",2010,7.9,"Centre-Est (FR)"
"Y_GE15","FR71",2010,8.1,"Rhône-Alpes"
"Y_GE15","FR72",2010,7,"Auvergne"
"Y_GE15","FR8",2010,10.9,"Méditerranée"
"Y_GE15","FR81",2010,13.7,"Languedoc-Roussillon"
"Y_GE15","FR82",2010,9.7,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2010,6,"Corse"
"Y_GE15","FRA",2010,25.2,"Départements d'outre-mer"
"Y_GE15","FRA1",2010,23.8,"Guadeloupe"
"Y_GE15","FRA2",2010,21,"Martinique"
"Y_GE15","FRA3",2010,21,"Guyane"
"Y_GE15","FRA4",2010,28.9,"La Réunion"
"Y_GE15","HR",2010,11.6,"Croatia"
"Y_GE15","HR0",2010,11.6,"Hrvatska"
"Y_GE15","HR03",2010,11.1,"Jadranska Hrvatska"
"Y_GE15","HR04",2010,11.9,"Kontinentalna Hrvatska"
"Y_GE15","HU",2010,11.2,"Hungary"
"Y_GE15","HU1",2010,8.9,"Közép-Magyarország"
"Y_GE15","HU10",2010,8.9,"Közép-Magyarország"
"Y_GE15","HU2",2010,10.5,"Dunántúl"
"Y_GE15","HU21",2010,10,"Közép-Dunántúl"
"Y_GE15","HU22",2010,9.3,"Nyugat-Dunántúl"
"Y_GE15","HU23",2010,12.4,"Dél-Dunántúl"
"Y_GE15","HU3",2010,13.6,"Alföld és Észak"
"Y_GE15","HU31",2010,16.2,"Észak-Magyarország"
"Y_GE15","HU32",2010,14.4,"Észak-Alföld"
"Y_GE15","HU33",2010,10.4,"Dél-Alföld"
"Y_GE15","IE",2010,13.9,"Ireland"
"Y_GE15","IE0",2010,13.9,"Éire/Ireland"
"Y_GE15","IE01",2010,14.5,"Border, Midland and Western"
"Y_GE15","IE02",2010,13.6,"Southern and Eastern"
"Y_GE15","IS",2010,7.6,"Iceland"
"Y_GE15","IS0",2010,7.6,"Ísland"
"Y_GE15","IS00",2010,7.6,"Ísland"
"Y_GE15","IT",2010,8.4,"Italy"
"Y_GE15","ITC",2010,6.2,"Nord-Ovest"
"Y_GE15","ITC1",2010,7.5,"Piemonte"
"Y_GE15","ITC2",2010,4.5,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2010,6.6,"Liguria"
"Y_GE15","ITC4",2010,5.5,"Lombardia"
"Y_GE15","ITF",2010,12.7,"Sud"
"Y_GE15","ITF1",2010,8.7,"Abruzzo"
"Y_GE15","ITF2",2010,8.4,"Molise"
"Y_GE15","ITF3",2010,13.9,"Campania"
"Y_GE15","ITF4",2010,13.5,"Puglia"
"Y_GE15","ITF5",2010,12.9,"Basilicata"
"Y_GE15","ITF6",2010,11.9,"Calabria"
"Y_GE15","ITG",2010,14.4,"Isole"
"Y_GE15","ITG1",2010,14.6,"Sicilia"
"Y_GE15","ITG2",2010,14,"Sardegna"
"Y_GE15","ITH",2010,5.4,"Nord-Est"
"Y_GE15","ITH1",2010,2.7,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2010,4.2,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2010,5.7,"Veneto"
"Y_GE15","ITH4",2010,5.7,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2010,5.6,"Emilia-Romagna"
"Y_GE15","ITI",2010,7.5,"Centro (IT)"
"Y_GE15","ITI1",2010,6,"Toscana"
"Y_GE15","ITI2",2010,6.6,"Umbria"
"Y_GE15","ITI3",2010,5.7,"Marche"
"Y_GE15","ITI4",2010,9.2,"Lazio"
"Y_GE15","LT",2010,17.8,"Lithuania"
"Y_GE15","LT0",2010,17.8,"Lietuva"
"Y_GE15","LT00",2010,17.8,"Lietuva"
"Y_GE15","LU",2010,4.4,"Luxembourg"
"Y_GE15","LU0",2010,4.4,"Luxembourg"
"Y_GE15","LU00",2010,4.4,"Luxembourg"
"Y_GE15","LV",2010,19.5,"Latvia"
"Y_GE15","LV0",2010,19.5,"Latvija"
"Y_GE15","LV00",2010,19.5,"Latvija"
"Y_GE15","MK",2010,32,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2010,32,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2010,32,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2010,6.8,"Malta"
"Y_GE15","MT0",2010,6.8,"Malta"
"Y_GE15","MT00",2010,6.8,"Malta"
"Y_GE15","NL",2010,4.5,"Netherlands"
"Y_GE15","NL1",2010,4.9,"Noord-Nederland"
"Y_GE15","NL11",2010,5.3,"Groningen"
"Y_GE15","NL12",2010,4.8,"Friesland (NL)"
"Y_GE15","NL13",2010,4.5,"Drenthe"
"Y_GE15","NL2",2010,4.3,"Oost-Nederland"
"Y_GE15","NL21",2010,4.4,"Overijssel"
"Y_GE15","NL22",2010,4.1,"Gelderland"
"Y_GE15","NL23",2010,5.2,"Flevoland"
"Y_GE15","NL3",2010,4.4,"West-Nederland"
"Y_GE15","NL31",2010,3.7,"Utrecht"
"Y_GE15","NL32",2010,4.2,"Noord-Holland"
"Y_GE15","NL33",2010,5,"Zuid-Holland"
"Y_GE15","NL34",2010,2.7,"Zeeland"
"Y_GE15","NL4",2010,4.5,"Zuid-Nederland"
"Y_GE15","NL41",2010,4.2,"Noord-Brabant"
"Y_GE15","NL42",2010,5.1,"Limburg (NL)"
"Y_GE15","NO",2010,3.5,"Norway"
"Y_GE15","NO0",2010,3.5,"Norge"
"Y_GE15","NO01",2010,4,"Oslo og Akershus"
"Y_GE15","NO02",2010,3.2,"Hedmark og Oppland"
"Y_GE15","NO03",2010,3.7,"Sør-Østlandet"
"Y_GE15","NO04",2010,2.6,"Agder og Rogaland"
"Y_GE15","NO05",2010,3.4,"Vestlandet"
"Y_GE15","NO06",2010,3.6,"Trøndelag"
"Y_GE15","NO07",2010,3.8,"Nord-Norge"
"Y_GE15","PL",2010,9.6,"Poland"
"Y_GE15","PL1",2010,8.1,"Region Centralny"
"Y_GE15","PL11",2010,9.3,"Lódzkie"
"Y_GE15","PL12",2010,7.4,"Mazowieckie"
"Y_GE15","PL2",2010,9.1,"Region Poludniowy"
"Y_GE15","PL21",2010,9.1,"Malopolskie"
"Y_GE15","PL22",2010,9.2,"Slaskie"
"Y_GE15","PL3",2010,10.9,"Region Wschodni"
"Y_GE15","PL31",2010,9.8,"Lubelskie"
"Y_GE15","PL32",2010,11.6,"Podkarpackie"
"Y_GE15","PL33",2010,12,"Swietokrzyskie"
"Y_GE15","PL34",2010,10.2,"Podlaskie"
"Y_GE15","PL4",2010,10,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2010,8.8,"Wielkopolskie"
"Y_GE15","PL42",2010,12.4,"Zachodniopomorskie"
"Y_GE15","PL43",2010,10.6,"Lubuskie"
"Y_GE15","PL5",2010,10.9,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2010,11.3,"Dolnoslaskie"
"Y_GE15","PL52",2010,9.6,"Opolskie"
"Y_GE15","PL6",2010,9.9,"Region Pólnocny"
"Y_GE15","PL61",2010,10.6,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2010,9.7,"Warminsko-Mazurskie"
"Y_GE15","PL63",2010,9.3,"Pomorskie"
"Y_GE15","PT",2010,10.8,"Portugal"
"Y_GE15","PT1",2010,10.9,"Continente"
"Y_GE15","PT11",2010,12.6,"Norte"
"Y_GE15","PT15",2010,13.4,"Algarve"
"Y_GE15","PT16",2010,7.6,"Centro (PT)"
"Y_GE15","PT17",2010,11.3,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2010,11.4,"Alentejo"
"Y_GE15","PT2",2010,6.8,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2010,6.8,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2010,7.4,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2010,7.4,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2010,7,"Romania"
"Y_GE15","RO1",2010,8.2,"Macroregiunea unu"
"Y_GE15","RO11",2010,6.5,"Nord-Vest"
"Y_GE15","RO12",2010,10.3,"Centru"
"Y_GE15","RO2",2010,6.6,"Macroregiunea doi"
"Y_GE15","RO21",2010,5.5,"Nord-Est"
"Y_GE15","RO22",2010,8.2,"Sud-Est"
"Y_GE15","RO3",2010,6.4,"Macroregiunea trei"
"Y_GE15","RO31",2010,7.8,"Sud - Muntenia"
"Y_GE15","RO32",2010,4.7,"Bucuresti - Ilfov"
"Y_GE15","RO4",2010,6.7,"Macroregiunea patru"
"Y_GE15","RO41",2010,7.3,"Sud-Vest Oltenia"
"Y_GE15","RO42",2010,6,"Vest"
"Y_GE15","SE",2010,8.6,"Sweden"
"Y_GE15","SE1",2010,8.2,"Östra Sverige"
"Y_GE15","SE11",2010,7.2,"Stockholm"
"Y_GE15","SE12",2010,9.7,"Östra Mellansverige"
"Y_GE15","SE2",2010,8.6,"Södra Sverige"
"Y_GE15","SE21",2010,7.9,"Småland med öarna"
"Y_GE15","SE22",2010,8.8,"Sydsverige"
"Y_GE15","SE23",2010,8.7,"Västsverige"
"Y_GE15","SE3",2010,9.4,"Norra Sverige"
"Y_GE15","SE31",2010,9,"Norra Mellansverige"
"Y_GE15","SE32",2010,10.3,"Mellersta Norrland"
"Y_GE15","SE33",2010,9.5,"Övre Norrland"
"Y_GE15","SI",2010,7.2,"Slovenia"
"Y_GE15","SI0",2010,7.2,"Slovenija"
"Y_GE15","SI03",2010,7.8,"Vzhodna Slovenija"
"Y_GE15","SI04",2010,6.6,"Zahodna Slovenija"
"Y_GE15","SK",2010,14.4,"Slovakia"
"Y_GE15","SK0",2010,14.4,"Slovensko"
"Y_GE15","SK01",2010,6.2,"Bratislavský kraj"
"Y_GE15","SK02",2010,12.7,"Západné Slovensko"
"Y_GE15","SK03",2010,16.5,"Stredné Slovensko"
"Y_GE15","SK04",2010,18.5,"Východné Slovensko"
"Y_GE15","TR",2010,10.7,"Turkey"
"Y_GE15","TR1",2010,13.5,"Istanbul"
"Y_GE15","TR10",2010,13.5,"Istanbul"
"Y_GE15","TR2",2010,7.3,"Bati Marmara"
"Y_GE15","TR21",2010,8.4,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2010,6,"Balikesir, Çanakkale"
"Y_GE15","TR3",2010,10.9,"Ege"
"Y_GE15","TR31",2010,14.1,"Izmir"
"Y_GE15","TR32",2010,10.3,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2010,6.8,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2010,10.1,"Dogu Marmara"
"Y_GE15","TR41",2010,9.2,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2010,11.1,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2010,9.5,"Bati Anadolu"
"Y_GE15","TR51",2010,10.7,"Ankara"
"Y_GE15","TR52",2010,7.1,"Konya, Karaman"
"Y_GE15","TR6",2010,12.4,"Akdeniz"
"Y_GE15","TR61",2010,9.8,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2010,14.9,"Adana, Mersin"
"Y_GE15","TR63",2010,11.7,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2010,10.9,"Orta Anadolu"
"Y_GE15","TR71",2010,9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2010,12.3,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2010,7.3,"Bati Karadeniz"
"Y_GE15","TR81",2010,10.2,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2010,7.5,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2010,6,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2010,4.8,"Dogu Karadeniz"
"Y_GE15","TR90",2010,4.8,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2010,7,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2010,5.5,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2010,8.7,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2010,12.9,"Ortadogu Anadolu"
"Y_GE15","TRB1",2010,10.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2010,15.5,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2010,11.1,"Güneydogu Anadolu"
"Y_GE15","TRC1",2010,11.4,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2010,11.1,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2010,10.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2010,7.8,"United Kingdom"
"Y_GE15","UKC",2010,9.4,"North East (UK)"
"Y_GE15","UKC1",2010,9.1,"Tees Valley and Durham"
"Y_GE15","UKC2",2010,9.6,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2010,7.9,"North West (UK)"
"Y_GE15","UKD1",2010,6.5,"Cumbria"
"Y_GE15","UKD3",2010,8.7,"Greater Manchester"
"Y_GE15","UKD4",2010,5.9,"Lancashire"
"Y_GE15","UKD6",2010,6.1,"Cheshire"
"Y_GE15","UKD7",2010,10.5,"Merseyside"
"Y_GE15","UKE",2010,9.1,"Yorkshire and The Humber"
"Y_GE15","UKE1",2010,9.4,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2010,6.7,"North Yorkshire"
"Y_GE15","UKE3",2010,9.4,"South Yorkshire"
"Y_GE15","UKE4",2010,9.7,"West Yorkshire"
"Y_GE15","UKF",2010,7.6,"East Midlands (UK)"
"Y_GE15","UKF1",2010,8.8,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2010,7.2,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2010,4.9,"Lincolnshire"
"Y_GE15","UKG",2010,9,"West Midlands (UK)"
"Y_GE15","UKG1",2010,6.3,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2010,7.7,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2010,11.1,"West Midlands"
"Y_GE15","UKH",2010,6.6,"East of England"
"Y_GE15","UKH1",2010,6.6,"East Anglia"
"Y_GE15","UKH2",2010,6,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2010,7,"Essex"
"Y_GE15","UKI",2010,9.2,"London"
"Y_GE15","UKI3",2010,8.1,"Inner London - West"
"Y_GE15","UKI4",2010,10.9,"Inner London - East"
"Y_GE15","UKI5",2010,10,"Outer London - East and North East"
"Y_GE15","UKI6",2010,7.1,"Outer London - South"
"Y_GE15","UKI7",2010,8.6,"Outer London - West and North West"
"Y_GE15","UKJ",2010,6.1,"South East (UK)"
"Y_GE15","UKJ1",2010,5.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2010,5.1,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2010,6.3,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2010,7.7,"Kent"
"Y_GE15","UKK",2010,5.9,"South West (UK)"
"Y_GE15","UKK1",2010,5.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2010,5.4,"Dorset and Somerset"
"Y_GE15","UKK3",2010,8.1,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2010,6.5,"Devon"
"Y_GE15","UKL",2010,8.6,"Wales"
"Y_GE15","UKL1",2010,9.2,"West Wales and The Valleys"
"Y_GE15","UKL2",2010,7.8,"East Wales"
"Y_GE15","UKM",2010,8.2,"Scotland"
"Y_GE15","UKM2",2010,7.8,"Eastern Scotland"
"Y_GE15","UKM3",2010,10.1,"South Western Scotland"
"Y_GE15","UKM5",2010,3.6,"North Eastern Scotland"
"Y_GE15","UKM6",2010,7,"Highlands and Islands"
"Y_GE15","UKN",2010,7.1,"Northern Ireland (UK)"
"Y_GE15","UKN0",2010,7.1,"Northern Ireland (UK)"
"Y_GE25","AT",2010,4.1,"Austria"
"Y_GE25","AT1",2010,5.1,"Ostösterreich"
"Y_GE25","AT11",2010,3.2,"Burgenland (AT)"
"Y_GE25","AT12",2010,3.4,"Niederösterreich"
"Y_GE25","AT13",2010,7.1,"Wien"
"Y_GE25","AT2",2010,3.7,"Südösterreich"
"Y_GE25","AT21",2010,3.7,"Kärnten"
"Y_GE25","AT22",2010,3.7,"Steiermark"
"Y_GE25","AT3",2010,3.1,"Westösterreich"
"Y_GE25","AT31",2010,3.3,"Oberösterreich"
"Y_GE25","AT32",2010,2.6,"Salzburg"
"Y_GE25","AT33",2010,2.6,"Tirol"
"Y_GE25","AT34",2010,3.6,"Vorarlberg"
"Y_GE25","BE",2010,6.9,"Belgium"
"Y_GE25","BE1",2010,15.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2010,15.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2010,4.2,"Vlaams Gewest"
"Y_GE25","BE21",2010,4.9,"Prov. Antwerpen"
"Y_GE25","BE22",2010,4.1,"Prov. Limburg (BE)"
"Y_GE25","BE23",2010,4.2,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2010,4.1,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2010,3.1,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2010,9.5,"Région wallonne"
"Y_GE25","BE31",2010,6.9,"Prov. Brabant Wallon"
"Y_GE25","BE32",2010,11.5,"Prov. Hainaut"
"Y_GE25","BE33",2010,9.9,"Prov. Liège"
"Y_GE25","BE34",2010,6,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2010,7.7,"Prov. Namur"
"Y_GE25","BG",2010,9.2,"Bulgaria"
"Y_GE25","BG3",2010,11,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2010,10.4,"Severozapaden"
"Y_GE25","BG32",2010,10.4,"Severen tsentralen"
"Y_GE25","BG33",2010,13.6,"Severoiztochen"
"Y_GE25","BG34",2010,9.5,"Yugoiztochen"
"Y_GE25","BG4",2010,7.6,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2010,6.1,"Yugozapaden"
"Y_GE25","BG42",2010,9.9,"Yuzhen tsentralen"
"Y_GE25","CH",2010,4,"Switzerland"
"Y_GE25","CH0",2010,4,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2010,5.7,"Région lémanique"
"Y_GE25","CH02",2010,3.7,"Espace Mittelland"
"Y_GE25","CH03",2010,3.9,"Nordwestschweiz"
"Y_GE25","CH04",2010,3.9,"Zürich"
"Y_GE25","CH05",2010,3.2,"Ostschweiz"
"Y_GE25","CH06",2010,2.7,"Zentralschweiz"
"Y_GE25","CH07",2010,5.5,"Ticino"
"Y_GE25","CY",2010,5.1,"Cyprus"
"Y_GE25","CY0",2010,5.1,"Kypros"
"Y_GE25","CY00",2010,5.1,"Kypros"
"Y_GE25","CZ",2010,6.4,"Czech Republic"
"Y_GE25","CZ0",2010,6.4,"Ceská republika"
"Y_GE25","CZ01",2010,3.4,"Praha"
"Y_GE25","CZ02",2010,4.3,"Strední Cechy"
"Y_GE25","CZ03",2010,4.7,"Jihozápad"
"Y_GE25","CZ04",2010,9.4,"Severozápad"
"Y_GE25","CZ05",2010,5.8,"Severovýchod"
"Y_GE25","CZ06",2010,6.7,"Jihovýchod"
"Y_GE25","CZ07",2010,7.9,"Strední Morava"
"Y_GE25","CZ08",2010,9.3,"Moravskoslezsko"
"Y_GE25","DE",2010,6.6,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2010,4.4,"Baden-Württemberg"
"Y_GE25","DE11",2010,4.7,"Stuttgart"
"Y_GE25","DE12",2010,4.8,"Karlsruhe"
"Y_GE25","DE13",2010,3.7,"Freiburg"
"Y_GE25","DE14",2010,4.3,"Tübingen"
"Y_GE25","DE2",2010,4,"Bayern"
"Y_GE25","DE21",2010,3.4,"Oberbayern"
"Y_GE25","DE22",2010,3.5,"Niederbayern"
"Y_GE25","DE23",2010,3.8,"Oberpfalz"
"Y_GE25","DE24",2010,5.5,"Oberfranken"
"Y_GE25","DE25",2010,5.1,"Mittelfranken"
"Y_GE25","DE26",2010,4.6,"Unterfranken"
"Y_GE25","DE27",2010,4,"Schwaben"
"Y_GE25","DE3",2010,12.4,"Berlin"
"Y_GE25","DE30",2010,12.4,"Berlin"
"Y_GE25","DE4",2010,9.3,"Brandenburg"
"Y_GE25","DE40",2010,9.3,"Brandenburg"
"Y_GE25","DE5",2010,7.9,"Bremen"
"Y_GE25","DE50",2010,7.9,"Bremen"
"Y_GE25","DE6",2010,7,"Hamburg"
"Y_GE25","DE60",2010,7,"Hamburg"
"Y_GE25","DE7",2010,5.2,"Hessen"
"Y_GE25","DE71",2010,5.3,"Darmstadt"
"Y_GE25","DE72",2010,5,"Gießen"
"Y_GE25","DE73",2010,5.3,"Kassel"
"Y_GE25","DE8",2010,12.2,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2010,12.2,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2010,5.9,"Niedersachsen"
"Y_GE25","DE91",2010,6.7,"Braunschweig"
"Y_GE25","DE92",2010,6.5,"Hannover"
"Y_GE25","DE93",2010,5.1,"Lüneburg"
"Y_GE25","DE94",2010,5.5,"Weser-Ems"
"Y_GE25","DEA",2010,6.9,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2010,7.1,"Düsseldorf"
"Y_GE25","DEA2",2010,6.6,"Köln"
"Y_GE25","DEA3",2010,6.3,"Münster"
"Y_GE25","DEA4",2010,6.6,"Detmold"
"Y_GE25","DEA5",2010,7.8,"Arnsberg"
"Y_GE25","DEB",2010,4.9,"Rheinland-Pfalz"
"Y_GE25","DEB1",2010,4.9,"Koblenz"
"Y_GE25","DEB2",2010,3.7,"Trier"
"Y_GE25","DEB3",2010,5.3,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2010,6.5,"Saarland"
"Y_GE25","DEC0",2010,6.5,"Saarland"
"Y_GE25","DED",2010,11,"Sachsen"
"Y_GE25","DED2",2010,10.1,"Dresden"
"Y_GE25","DED4",2010,11.4,"Chemnitz"
"Y_GE25","DED5",2010,11.8,"Leipzig"
"Y_GE25","DEE",2010,11.2,"Sachsen-Anhalt"
"Y_GE25","DEE0",2010,11.2,"Sachsen-Anhalt"
"Y_GE25","DEF",2010,6.2,"Schleswig-Holstein"
"Y_GE25","DEF0",2010,6.2,"Schleswig-Holstein"
"Y_GE25","DEG",2010,8.4,"Thüringen"
"Y_GE25","DEG0",2010,8.4,"Thüringen"
"Y_GE25","DK",2010,6.3,"Denmark"
"Y_GE25","DK0",2010,6.3,"Danmark"
"Y_GE25","DK01",2010,6.7,"Hovedstaden"
"Y_GE25","DK02",2010,5.3,"Sjælland"
"Y_GE25","DK03",2010,6.3,"Syddanmark"
"Y_GE25","DK04",2010,6,"Midtjylland"
"Y_GE25","DK05",2010,6.7,"Nordjylland"
"Y_GE25","EA17",2010,8.8,"Euro area (17 countries)"
"Y_GE25","EA18",2010,8.9,"Euro area (18 countries)"
"Y_GE25","EA19",2010,8.9,"Euro area (19 countries)"
"Y_GE25","EE",2010,14.9,"Estonia"
"Y_GE25","EE0",2010,14.9,"Eesti"
"Y_GE25","EE00",2010,14.9,"Eesti"
"Y_GE25","EL",2010,11.2,"Greece"
"Y_GE25","EL3",2010,11.3,"Attiki"
"Y_GE25","EL30",2010,11.3,"Attiki"
"Y_GE25","EL4",2010,10.7,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2010,7.6,"Voreio Aigaio"
"Y_GE25","EL42",2010,13.1,"Notio Aigaio"
"Y_GE25","EL43",2010,10.4,"Kriti"
"Y_GE25","EL5",2010,12.3,"Voreia Ellada"
"Y_GE25","EL51",2010,12.3,"Anatoliki Makedonia, Thraki"
"Y_GE25","EL52",2010,12.3,"Kentriki Makedonia"
"Y_GE25","EL53",2010,14.3,"Dytiki Makedonia"
"Y_GE25","EL54",2010,10.6,"Ipeiros"
"Y_GE25","EL6",2010,9.9,"Kentriki Ellada"
"Y_GE25","EL61",2010,10.1,"Thessalia"
"Y_GE25","EL62",2010,12.9,"Ionia Nisia"
"Y_GE25","EL63",2010,9.7,"Dytiki Ellada"
"Y_GE25","EL64",2010,10.4,"Sterea Ellada"
"Y_GE25","EL65",2010,8.4,"Peloponnisos"
"Y_GE25","ES",2010,17.8,"Spain"
"Y_GE25","ES1",2010,13.7,"Noroeste (ES)"
"Y_GE25","ES11",2010,13.8,"Galicia"
"Y_GE25","ES12",2010,14.5,"Principado de Asturias"
"Y_GE25","ES13",2010,12,"Cantabria"
"Y_GE25","ES2",2010,10.9,"Noreste (ES)"
"Y_GE25","ES21",2010,9.4,"País Vasco"
"Y_GE25","ES22",2010,10.3,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2010,12.4,"La Rioja"
"Y_GE25","ES24",2010,13.5,"Aragón"
"Y_GE25","ES3",2010,14,"Comunidad de Madrid"
"Y_GE25","ES30",2010,14,"Comunidad de Madrid"
"Y_GE25","ES4",2010,16.9,"Centro (ES)"
"Y_GE25","ES41",2010,14.2,"Castilla y León"
"Y_GE25","ES42",2010,18.6,"Castilla-la Mancha"
"Y_GE25","ES43",2010,20.2,"Extremadura"
"Y_GE25","ES5",2010,17.6,"Este (ES)"
"Y_GE25","ES51",2010,15.6,"Cataluña"
"Y_GE25","ES52",2010,20.9,"Comunidad Valenciana"
"Y_GE25","ES53",2010,17.8,"Illes Balears"
"Y_GE25","ES6",2010,24.4,"Sur (ES)"
"Y_GE25","ES61",2010,25.2,"Andalucía"
"Y_GE25","ES62",2010,21,"Región de Murcia"
"Y_GE25","ES63",2010,19,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2010,19,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2010,26.3,"Canarias (ES)"
"Y_GE25","ES70",2010,26.3,"Canarias (ES)"
"Y_GE25","EU15",2010,8.2,"European Union (15 countries)"
"Y_GE25","EU27",2010,8.2,"European Union (27 countries)"
"Y_GE25","EU28",2010,8.2,"European Union (28 countries)"
"Y_GE25","FI",2010,6.6,"Finland"
"Y_GE25","FI1",2010,6.7,"Manner-Suomi"
"Y_GE25","FI19",2010,7,"Länsi-Suomi"
"Y_GE25","FI1B",2010,4.7,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2010,7.5,"Etelä-Suomi"
"Y_GE25","FI1D",2010,8.2,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2010,NA,"Åland"
"Y_GE25","FI20",2010,NA,"Åland"
"Y_GE25","FR",2010,7.7,"France"
"Y_GE25","FR1",2010,7.4,"Île de France"
"Y_GE25","FR10",2010,7.4,"Île de France"
"Y_GE25","FR2",2010,7.2,"Bassin Parisien"
"Y_GE25","FR21",2010,7,"Champagne-Ardenne"
"Y_GE25","FR22",2010,9.3,"Picardie"
"Y_GE25","FR23",2010,7.4,"Haute-Normandie"
"Y_GE25","FR24",2010,5.9,"Centre (FR)"
"Y_GE25","FR25",2010,6.7,"Basse-Normandie"
"Y_GE25","FR26",2010,7.3,"Bourgogne"
"Y_GE25","FR3",2010,10.2,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2010,10.2,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2010,6.9,"Est (FR)"
"Y_GE25","FR41",2010,7.3,"Lorraine"
"Y_GE25","FR42",2010,6.7,"Alsace"
"Y_GE25","FR43",2010,6.8,"Franche-Comté"
"Y_GE25","FR5",2010,6.4,"Ouest (FR)"
"Y_GE25","FR51",2010,7.2,"Pays de la Loire"
"Y_GE25","FR52",2010,5.6,"Bretagne"
"Y_GE25","FR53",2010,6.4,"Poitou-Charentes"
"Y_GE25","FR6",2010,6.4,"Sud-Ouest (FR)"
"Y_GE25","FR61",2010,6.5,"Aquitaine"
"Y_GE25","FR62",2010,6.3,"Midi-Pyrénées"
"Y_GE25","FR63",2010,5.8,"Limousin"
"Y_GE25","FR7",2010,6.4,"Centre-Est (FR)"
"Y_GE25","FR71",2010,6.6,"Rhône-Alpes"
"Y_GE25","FR72",2010,5.4,"Auvergne"
"Y_GE25","FR8",2010,9,"Méditerranée"
"Y_GE25","FR81",2010,11.3,"Languedoc-Roussillon"
"Y_GE25","FR82",2010,8,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2010,5.8,"Corse"
"Y_GE25","FRA",2010,21.5,"Départements d'outre-mer"
"Y_GE25","FRA1",2010,21.2,"Guadeloupe"
"Y_GE25","FRA2",2010,17.4,"Martinique"
"Y_GE25","FRA3",2010,18,"Guyane"
"Y_GE25","FRA4",2010,24.7,"La Réunion"
"Y_GE25","HR",2010,9.4,"Croatia"
"Y_GE25","HR0",2010,9.4,"Hrvatska"
"Y_GE25","HR03",2010,9.4,"Jadranska Hrvatska"
"Y_GE25","HR04",2010,9.4,"Kontinentalna Hrvatska"
"Y_GE25","HU",2010,10,"Hungary"
"Y_GE25","HU1",2010,8.2,"Közép-Magyarország"
"Y_GE25","HU10",2010,8.2,"Közép-Magyarország"
"Y_GE25","HU2",2010,9.3,"Dunántúl"
"Y_GE25","HU21",2010,9,"Közép-Dunántúl"
"Y_GE25","HU22",2010,8.2,"Nyugat-Dunántúl"
"Y_GE25","HU23",2010,11.1,"Dél-Dunántúl"
"Y_GE25","HU3",2010,12.1,"Alföld és Észak"
"Y_GE25","HU31",2010,14.9,"Észak-Magyarország"
"Y_GE25","HU32",2010,12.5,"Észak-Alföld"
"Y_GE25","HU33",2010,9.3,"Dél-Alföld"
"Y_GE25","IE",2010,12,"Ireland"
"Y_GE25","IE0",2010,12,"Éire/Ireland"
"Y_GE25","IE01",2010,12.4,"Border, Midland and Western"
"Y_GE25","IE02",2010,11.8,"Southern and Eastern"
"Y_GE25","IS",2010,5.8,"Iceland"
"Y_GE25","IS0",2010,5.8,"Ísland"
"Y_GE25","IS00",2010,5.8,"Ísland"
"Y_GE25","IT",2010,6.9,"Italy"
"Y_GE25","ITC",2010,5.1,"Nord-Ovest"
"Y_GE25","ITC1",2010,6.2,"Piemonte"
"Y_GE25","ITC2",2010,3.6,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2010,5.8,"Liguria"
"Y_GE25","ITC4",2010,4.6,"Lombardia"
"Y_GE25","ITF",2010,10.5,"Sud"
"Y_GE25","ITF1",2010,7.4,"Abruzzo"
"Y_GE25","ITF2",2010,6.8,"Molise"
"Y_GE25","ITF3",2010,11.3,"Campania"
"Y_GE25","ITF4",2010,11.2,"Puglia"
"Y_GE25","ITF5",2010,10.8,"Basilicata"
"Y_GE25","ITF6",2010,9.9,"Calabria"
"Y_GE25","ITG",2010,12,"Isole"
"Y_GE25","ITG1",2010,12,"Sicilia"
"Y_GE25","ITG2",2010,11.9,"Sardegna"
"Y_GE25","ITH",2010,4.5,"Nord-Est"
"Y_GE25","ITH1",2010,2.3,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2010,3.4,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2010,4.7,"Veneto"
"Y_GE25","ITH4",2010,5,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2010,4.6,"Emilia-Romagna"
"Y_GE25","ITI",2010,6.4,"Centro (IT)"
"Y_GE25","ITI1",2010,5,"Toscana"
"Y_GE25","ITI2",2010,5.6,"Umbria"
"Y_GE25","ITI3",2010,5,"Marche"
"Y_GE25","ITI4",2010,7.8,"Lazio"
"Y_GE25","LT",2010,16.1,"Lithuania"
"Y_GE25","LT0",2010,16.1,"Lietuva"
"Y_GE25","LT00",2010,16.1,"Lietuva"
"Y_GE25","LU",2010,3.7,"Luxembourg"
"Y_GE25","LU0",2010,3.7,"Luxembourg"
"Y_GE25","LU00",2010,3.7,"Luxembourg"
"Y_GE25","LV",2010,17.4,"Latvia"
"Y_GE25","LV0",2010,17.4,"Latvija"
"Y_GE25","LV00",2010,17.4,"Latvija"
"Y_GE25","MK",2010,29.3,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2010,29.3,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2010,29.3,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2010,5.6,"Malta"
"Y_GE25","MT0",2010,5.6,"Malta"
"Y_GE25","MT00",2010,5.6,"Malta"
"Y_GE25","NL",2010,3.7,"Netherlands"
"Y_GE25","NL1",2010,4,"Noord-Nederland"
"Y_GE25","NL11",2010,4.3,"Groningen"
"Y_GE25","NL12",2010,4,"Friesland (NL)"
"Y_GE25","NL13",2010,3.7,"Drenthe"
"Y_GE25","NL2",2010,3.4,"Oost-Nederland"
"Y_GE25","NL21",2010,3.6,"Overijssel"
"Y_GE25","NL22",2010,3.3,"Gelderland"
"Y_GE25","NL23",2010,3.8,"Flevoland"
"Y_GE25","NL3",2010,3.6,"West-Nederland"
"Y_GE25","NL31",2010,3,"Utrecht"
"Y_GE25","NL32",2010,3.5,"Noord-Holland"
"Y_GE25","NL33",2010,4.1,"Zuid-Holland"
"Y_GE25","NL34",2010,2.5,"Zeeland"
"Y_GE25","NL4",2010,3.8,"Zuid-Nederland"
"Y_GE25","NL41",2010,3.6,"Noord-Brabant"
"Y_GE25","NL42",2010,4.3,"Limburg (NL)"
"Y_GE25","NO",2010,2.6,"Norway"
"Y_GE25","NO0",2010,2.6,"Norge"
"Y_GE25","NO01",2010,3.2,"Oslo og Akershus"
"Y_GE25","NO02",2010,2,"Hedmark og Oppland"
"Y_GE25","NO03",2010,2.7,"Sør-Østlandet"
"Y_GE25","NO04",2010,2.1,"Agder og Rogaland"
"Y_GE25","NO05",2010,2.5,"Vestlandet"
"Y_GE25","NO06",2010,2.4,"Trøndelag"
"Y_GE25","NO07",2010,2.4,"Nord-Norge"
"Y_GE25","PL",2010,8,"Poland"
"Y_GE25","PL1",2010,6.9,"Region Centralny"
"Y_GE25","PL11",2010,8,"Lódzkie"
"Y_GE25","PL12",2010,6.3,"Mazowieckie"
"Y_GE25","PL2",2010,7.6,"Region Poludniowy"
"Y_GE25","PL21",2010,7.5,"Malopolskie"
"Y_GE25","PL22",2010,7.6,"Slaskie"
"Y_GE25","PL3",2010,8.9,"Region Wschodni"
"Y_GE25","PL31",2010,8.3,"Lubelskie"
"Y_GE25","PL32",2010,9,"Podkarpackie"
"Y_GE25","PL33",2010,10.2,"Swietokrzyskie"
"Y_GE25","PL34",2010,8.6,"Podlaskie"
"Y_GE25","PL4",2010,8.3,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2010,6.9,"Wielkopolskie"
"Y_GE25","PL42",2010,10.6,"Zachodniopomorskie"
"Y_GE25","PL43",2010,9.1,"Lubuskie"
"Y_GE25","PL5",2010,9.4,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2010,9.8,"Dolnoslaskie"
"Y_GE25","PL52",2010,8.1,"Opolskie"
"Y_GE25","PL6",2010,8.3,"Region Pólnocny"
"Y_GE25","PL61",2010,8.7,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2010,8.2,"Warminsko-Mazurskie"
"Y_GE25","PL63",2010,7.9,"Pomorskie"
"Y_GE25","PT",2010,9.8,"Portugal"
"Y_GE25","PT1",2010,10,"Continente"
"Y_GE25","PT11",2010,11.6,"Norte"
"Y_GE25","PT15",2010,12.1,"Algarve"
"Y_GE25","PT16",2010,6.9,"Centro (PT)"
"Y_GE25","PT17",2010,10.3,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2010,10.1,"Alentejo"
"Y_GE25","PT2",2010,5.4,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2010,5.4,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2010,6.4,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2010,6.4,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2010,5.6,"Romania"
"Y_GE25","RO1",2010,6.6,"Macroregiunea unu"
"Y_GE25","RO11",2010,5.3,"Nord-Vest"
"Y_GE25","RO12",2010,8.2,"Centru"
"Y_GE25","RO2",2010,5.4,"Macroregiunea doi"
"Y_GE25","RO21",2010,4.6,"Nord-Est"
"Y_GE25","RO22",2010,6.6,"Sud-Est"
"Y_GE25","RO3",2010,4.8,"Macroregiunea trei"
"Y_GE25","RO31",2010,5.7,"Sud - Muntenia"
"Y_GE25","RO32",2010,3.5,"Bucuresti - Ilfov"
"Y_GE25","RO4",2010,5.7,"Macroregiunea patru"
"Y_GE25","RO41",2010,6.4,"Sud-Vest Oltenia"
"Y_GE25","RO42",2010,4.9,"Vest"
"Y_GE25","SE",2010,6.2,"Sweden"
"Y_GE25","SE1",2010,6.1,"Östra Sverige"
"Y_GE25","SE11",2010,5.4,"Stockholm"
"Y_GE25","SE12",2010,7.1,"Östra Mellansverige"
"Y_GE25","SE2",2010,6.1,"Södra Sverige"
"Y_GE25","SE21",2010,5.7,"Småland med öarna"
"Y_GE25","SE22",2010,6.2,"Sydsverige"
"Y_GE25","SE23",2010,6.2,"Västsverige"
"Y_GE25","SE3",2010,6.7,"Norra Sverige"
"Y_GE25","SE31",2010,6.5,"Norra Mellansverige"
"Y_GE25","SE32",2010,7,"Mellersta Norrland"
"Y_GE25","SE33",2010,6.8,"Övre Norrland"
"Y_GE25","SI",2010,6.5,"Slovenia"
"Y_GE25","SI0",2010,6.5,"Slovenija"
"Y_GE25","SI03",2010,7.1,"Vzhodna Slovenija"
"Y_GE25","SI04",2010,5.8,"Zahodna Slovenija"
"Y_GE25","SK",2010,12.5,"Slovakia"
"Y_GE25","SK0",2010,12.5,"Slovensko"
"Y_GE25","SK01",2010,5.5,"Bratislavský kraj"
"Y_GE25","SK02",2010,10.9,"Západné Slovensko"
"Y_GE25","SK03",2010,14.4,"Stredné Slovensko"
"Y_GE25","SK04",2010,16.1,"Východné Slovensko"
"Y_GE25","TR",2010,8.8,"Turkey"
"Y_GE25","TR1",2010,11.6,"Istanbul"
"Y_GE25","TR10",2010,11.6,"Istanbul"
"Y_GE25","TR2",2010,6,"Bati Marmara"
"Y_GE25","TR21",2010,6.7,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2010,5.1,"Balikesir, Çanakkale"
"Y_GE25","TR3",2010,8.8,"Ege"
"Y_GE25","TR31",2010,11.6,"Izmir"
"Y_GE25","TR32",2010,8.4,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2010,5.1,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2010,8.3,"Dogu Marmara"
"Y_GE25","TR41",2010,7.6,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2010,9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2010,7.7,"Bati Anadolu"
"Y_GE25","TR51",2010,8.7,"Ankara"
"Y_GE25","TR52",2010,5.6,"Konya, Karaman"
"Y_GE25","TR6",2010,10.4,"Akdeniz"
"Y_GE25","TR61",2010,8,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2010,12.6,"Adana, Mersin"
"Y_GE25","TR63",2010,10,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2010,9,"Orta Anadolu"
"Y_GE25","TR71",2010,7.4,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2010,10.1,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2010,5.9,"Bati Karadeniz"
"Y_GE25","TR81",2010,7.4,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2010,6.1,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2010,5.2,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2010,3.5,"Dogu Karadeniz"
"Y_GE25","TR90",2010,3.5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2010,5.5,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2010,4.1,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2010,7.2,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2010,10,"Ortadogu Anadolu"
"Y_GE25","TRB1",2010,8.2,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2010,12.2,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2010,9.7,"Güneydogu Anadolu"
"Y_GE25","TRC1",2010,9.9,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2010,10.3,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2010,8.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2010,5.7,"United Kingdom"
"Y_GE25","UKC",2010,7.2,"North East (UK)"
"Y_GE25","UKC1",2010,7,"Tees Valley and Durham"
"Y_GE25","UKC2",2010,7.4,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2010,5.6,"North West (UK)"
"Y_GE25","UKD1",2010,3.8,"Cumbria"
"Y_GE25","UKD3",2010,6,"Greater Manchester"
"Y_GE25","UKD4",2010,4.2,"Lancashire"
"Y_GE25","UKD6",2010,4.4,"Cheshire"
"Y_GE25","UKD7",2010,7.9,"Merseyside"
"Y_GE25","UKE",2010,6.9,"Yorkshire and The Humber"
"Y_GE25","UKE1",2010,6.7,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2010,4.9,"North Yorkshire"
"Y_GE25","UKE3",2010,7.6,"South Yorkshire"
"Y_GE25","UKE4",2010,7.3,"West Yorkshire"
"Y_GE25","UKF",2010,5.7,"East Midlands (UK)"
"Y_GE25","UKF1",2010,6.7,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2010,5.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2010,3.8,"Lincolnshire"
"Y_GE25","UKG",2010,6.6,"West Midlands (UK)"
"Y_GE25","UKG1",2010,3.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2010,6.1,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2010,8.4,"West Midlands"
"Y_GE25","UKH",2010,4.9,"East of England"
"Y_GE25","UKH1",2010,4.7,"East Anglia"
"Y_GE25","UKH2",2010,4.4,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2010,5.6,"Essex"
"Y_GE25","UKI",2010,7.1,"London"
"Y_GE25","UKI3",2010,6.7,"Inner London - West"
"Y_GE25","UKI4",2010,8.1,"Inner London - East"
"Y_GE25","UKI5",2010,7.4,"Outer London - East and North East"
"Y_GE25","UKI6",2010,5.6,"Outer London - South"
"Y_GE25","UKI7",2010,6.9,"Outer London - West and North West"
"Y_GE25","UKJ",2010,4.5,"South East (UK)"
"Y_GE25","UKJ1",2010,4.7,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2010,3.9,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2010,4.5,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2010,5.1,"Kent"
"Y_GE25","UKK",2010,4.3,"South West (UK)"
"Y_GE25","UKK1",2010,3.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2010,4.3,"Dorset and Somerset"
"Y_GE25","UKK3",2010,5.5,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2010,4.5,"Devon"
"Y_GE25","UKL",2010,5.7,"Wales"
"Y_GE25","UKL1",2010,5.9,"West Wales and The Valleys"
"Y_GE25","UKL2",2010,5.5,"East Wales"
"Y_GE25","UKM",2010,6.1,"Scotland"
"Y_GE25","UKM2",2010,5.4,"Eastern Scotland"
"Y_GE25","UKM3",2010,7.9,"South Western Scotland"
"Y_GE25","UKM5",2010,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2010,5.3,"Highlands and Islands"
"Y_GE25","UKN",2010,5.1,"Northern Ireland (UK)"
"Y_GE25","UKN0",2010,5.1,"Northern Ireland (UK)"
"Y15-24","AT",2009,10.7,"Austria"
"Y15-24","AT1",2009,13.7,"Ostösterreich"
"Y15-24","AT11",2009,NA,"Burgenland (AT)"
"Y15-24","AT12",2009,12,"Niederösterreich"
"Y15-24","AT13",2009,16.3,"Wien"
"Y15-24","AT2",2009,10.4,"Südösterreich"
"Y15-24","AT21",2009,9.8,"Kärnten"
"Y15-24","AT22",2009,10.7,"Steiermark"
"Y15-24","AT3",2009,8,"Westösterreich"
"Y15-24","AT31",2009,7.6,"Oberösterreich"
"Y15-24","AT32",2009,8.1,"Salzburg"
"Y15-24","AT33",2009,6.9,"Tirol"
"Y15-24","AT34",2009,11.6,"Vorarlberg"
"Y15-24","BE",2009,21.9,"Belgium"
"Y15-24","BE1",2009,31.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2009,31.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2009,15.7,"Vlaams Gewest"
"Y15-24","BE21",2009,16.2,"Prov. Antwerpen"
"Y15-24","BE22",2009,18,"Prov. Limburg (BE)"
"Y15-24","BE23",2009,13.9,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2009,18.7,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2009,13,"Prov. West-Vlaanderen"
"Y15-24","BE3",2009,30.5,"Région wallonne"
"Y15-24","BE31",2009,19.4,"Prov. Brabant Wallon"
"Y15-24","BE32",2009,38,"Prov. Hainaut"
"Y15-24","BE33",2009,29.7,"Prov. Liège"
"Y15-24","BE34",2009,21.7,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2009,22.7,"Prov. Namur"
"Y15-24","BG",2009,16.2,"Bulgaria"
"Y15-24","BG3",2009,19.8,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2009,15.1,"Severozapaden"
"Y15-24","BG32",2009,21.7,"Severen tsentralen"
"Y15-24","BG33",2009,23.5,"Severoiztochen"
"Y15-24","BG34",2009,18,"Yugoiztochen"
"Y15-24","BG4",2009,12.7,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2009,10,"Yugozapaden"
"Y15-24","BG42",2009,17.3,"Yuzhen tsentralen"
"Y15-24","CH",2009,8.5,"Switzerland"
"Y15-24","CH0",2009,8.5,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2009,13.6,"Région lémanique"
"Y15-24","CH02",2009,8.3,"Espace Mittelland"
"Y15-24","CH03",2009,8.8,"Nordwestschweiz"
"Y15-24","CH04",2009,7.8,"Zürich"
"Y15-24","CH05",2009,4.6,"Ostschweiz"
"Y15-24","CH06",2009,5.4,"Zentralschweiz"
"Y15-24","CH07",2009,14.3,"Ticino"
"Y15-24","CY",2009,13.8,"Cyprus"
"Y15-24","CY0",2009,13.8,"Kypros"
"Y15-24","CY00",2009,13.8,"Kypros"
"Y15-24","CZ",2009,16.6,"Czech Republic"
"Y15-24","CZ0",2009,16.6,"Ceská republika"
"Y15-24","CZ01",2009,9.4,"Praha"
"Y15-24","CZ02",2009,15.3,"Strední Cechy"
"Y15-24","CZ03",2009,13.5,"Jihozápad"
"Y15-24","CZ04",2009,23.5,"Severozápad"
"Y15-24","CZ05",2009,14.9,"Severovýchod"
"Y15-24","CZ06",2009,15.8,"Jihovýchod"
"Y15-24","CZ07",2009,18.1,"Strední Morava"
"Y15-24","CZ08",2009,21.3,"Moravskoslezsko"
"Y15-24","DE",2009,11.2,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2009,8.3,"Baden-Württemberg"
"Y15-24","DE11",2009,9.5,"Stuttgart"
"Y15-24","DE12",2009,9.8,"Karlsruhe"
"Y15-24","DE13",2009,6.7,"Freiburg"
"Y15-24","DE14",2009,5.8,"Tübingen"
"Y15-24","DE2",2009,8.1,"Bayern"
"Y15-24","DE21",2009,6.4,"Oberbayern"
"Y15-24","DE22",2009,7.3,"Niederbayern"
"Y15-24","DE23",2009,7,"Oberpfalz"
"Y15-24","DE24",2009,13.6,"Oberfranken"
"Y15-24","DE25",2009,9.4,"Mittelfranken"
"Y15-24","DE26",2009,9.7,"Unterfranken"
"Y15-24","DE27",2009,7.1,"Schwaben"
"Y15-24","DE3",2009,17.5,"Berlin"
"Y15-24","DE30",2009,17.5,"Berlin"
"Y15-24","DE4",2009,17.2,"Brandenburg"
"Y15-24","DE40",2009,17.2,"Brandenburg"
"Y15-24","DE5",2009,NA,"Bremen"
"Y15-24","DE50",2009,NA,"Bremen"
"Y15-24","DE6",2009,10.4,"Hamburg"
"Y15-24","DE60",2009,10.4,"Hamburg"
"Y15-24","DE7",2009,11.3,"Hessen"
"Y15-24","DE71",2009,10.8,"Darmstadt"
"Y15-24","DE72",2009,12.9,"Gießen"
"Y15-24","DE73",2009,11.3,"Kassel"
"Y15-24","DE8",2009,15.1,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2009,15.1,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2009,10.3,"Niedersachsen"
"Y15-24","DE91",2009,10.8,"Braunschweig"
"Y15-24","DE92",2009,11.9,"Hannover"
"Y15-24","DE93",2009,9.5,"Lüneburg"
"Y15-24","DE94",2009,9.3,"Weser-Ems"
"Y15-24","DEA",2009,12.3,"Nordrhein-Westfalen"
"Y15-24","DEA1",2009,13.1,"Düsseldorf"
"Y15-24","DEA2",2009,10.6,"Köln"
"Y15-24","DEA3",2009,10.8,"Münster"
"Y15-24","DEA4",2009,12.1,"Detmold"
"Y15-24","DEA5",2009,14.1,"Arnsberg"
"Y15-24","DEB",2009,10.8,"Rheinland-Pfalz"
"Y15-24","DEB1",2009,10.9,"Koblenz"
"Y15-24","DEB2",2009,NA,"Trier"
"Y15-24","DEB3",2009,11.7,"Rheinhessen-Pfalz"
"Y15-24","DEC",2009,14.8,"Saarland"
"Y15-24","DEC0",2009,14.8,"Saarland"
"Y15-24","DED",2009,15,"Sachsen"
"Y15-24","DED2",2009,16.5,"Dresden"
"Y15-24","DED4",2009,13.2,"Chemnitz"
"Y15-24","DED5",2009,14.9,"Leipzig"
"Y15-24","DEE",2009,16.1,"Sachsen-Anhalt"
"Y15-24","DEE0",2009,16.1,"Sachsen-Anhalt"
"Y15-24","DEF",2009,10.6,"Schleswig-Holstein"
"Y15-24","DEF0",2009,10.6,"Schleswig-Holstein"
"Y15-24","DEG",2009,11.5,"Thüringen"
"Y15-24","DEG0",2009,11.5,"Thüringen"
"Y15-24","DK",2009,11.8,"Denmark"
"Y15-24","DK0",2009,11.8,"Danmark"
"Y15-24","DK01",2009,12.2,"Hovedstaden"
"Y15-24","DK02",2009,12.1,"Sjælland"
"Y15-24","DK03",2009,12,"Syddanmark"
"Y15-24","DK04",2009,11.2,"Midtjylland"
"Y15-24","DK05",2009,11.4,"Nordjylland"
"Y15-24","EA17",2009,20,"Euro area (17 countries)"
"Y15-24","EA18",2009,20.1,"Euro area (18 countries)"
"Y15-24","EA19",2009,20.1,"Euro area (19 countries)"
"Y15-24","EE",2009,27.4,"Estonia"
"Y15-24","EE0",2009,27.4,"Eesti"
"Y15-24","EE00",2009,27.4,"Eesti"
"Y15-24","EL",2009,25.7,"Greece"
"Y15-24","EL1",2009,28.6,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2009,30.4,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2009,28,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2009,34.8,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2009,26.6,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2009,29.8,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2009,34.7,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2009,26.5,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2009,28.8,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2009,32.9,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2009,25.8,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2009,21.9,"Attiki"
"Y15-24","EL30",2009,21.9,"Attiki"
"Y15-24","EL4",2009,22.5,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2009,24.6,"Voreio Aigaio"
"Y15-24","EL42",2009,24.5,"Notio Aigaio"
"Y15-24","EL43",2009,20.9,"Kriti"
"Y15-24","ES",2009,37.7,"Spain"
"Y15-24","ES1",2009,31.4,"Noroeste (ES)"
"Y15-24","ES11",2009,30.4,"Galicia"
"Y15-24","ES12",2009,35,"Principado de Asturias"
"Y15-24","ES13",2009,30,"Cantabria"
"Y15-24","ES2",2009,31.6,"Noreste (ES)"
"Y15-24","ES21",2009,31.6,"País Vasco"
"Y15-24","ES22",2009,30.6,"Comunidad Foral de Navarra"
"Y15-24","ES23",2009,33.1,"La Rioja"
"Y15-24","ES24",2009,31.7,"Aragón"
"Y15-24","ES3",2009,34.2,"Comunidad de Madrid"
"Y15-24","ES30",2009,34.2,"Comunidad de Madrid"
"Y15-24","ES4",2009,35.7,"Centro (ES)"
"Y15-24","ES41",2009,32,"Castilla y León"
"Y15-24","ES42",2009,36.3,"Castilla-la Mancha"
"Y15-24","ES43",2009,41.4,"Extremadura"
"Y15-24","ES5",2009,37.5,"Este (ES)"
"Y15-24","ES51",2009,36.9,"Cataluña"
"Y15-24","ES52",2009,39.5,"Comunidad Valenciana"
"Y15-24","ES53",2009,32.1,"Illes Balears"
"Y15-24","ES6",2009,43.3,"Sur (ES)"
"Y15-24","ES61",2009,45,"Andalucía"
"Y15-24","ES62",2009,33.7,"Región de Murcia"
"Y15-24","ES63",2009,35.7,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2009,38.3,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2009,47.8,"Canarias (ES)"
"Y15-24","ES70",2009,47.8,"Canarias (ES)"
"Y15-24","EU15",2009,19.7,"European Union (15 countries)"
"Y15-24","EU27",2009,20,"European Union (27 countries)"
"Y15-24","EU28",2009,20,"European Union (28 countries)"
"Y15-24","FI",2009,21.5,"Finland"
"Y15-24","FI1",2009,21.5,"Manner-Suomi"
"Y15-24","FI19",2009,21.7,"Länsi-Suomi"
"Y15-24","FI1B",2009,18.3,"Helsinki-Uusimaa"
"Y15-24","FI1C",2009,22.5,"Etelä-Suomi"
"Y15-24","FI1D",2009,24.7,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2009,NA,"Åland"
"Y15-24","FI20",2009,NA,"Åland"
"Y15-24","FR",2009,23.7,"France"
"Y15-24","FR1",2009,19.8,"Île de France"
"Y15-24","FR10",2009,19.8,"Île de France"
"Y15-24","FR2",2009,23.1,"Bassin Parisien"
"Y15-24","FR21",2009,20.3,"Champagne-Ardenne"
"Y15-24","FR22",2009,28.4,"Picardie"
"Y15-24","FR23",2009,23.9,"Haute-Normandie"
"Y15-24","FR24",2009,18.9,"Centre (FR)"
"Y15-24","FR25",2009,21.6,"Basse-Normandie"
"Y15-24","FR26",2009,26.9,"Bourgogne"
"Y15-24","FR3",2009,36.7,"Nord - Pas-de-Calais"
"Y15-24","FR30",2009,36.7,"Nord - Pas-de-Calais"
"Y15-24","FR4",2009,23.3,"Est (FR)"
"Y15-24","FR41",2009,27.5,"Lorraine"
"Y15-24","FR42",2009,20.1,"Alsace"
"Y15-24","FR43",2009,19.8,"Franche-Comté"
"Y15-24","FR5",2009,19,"Ouest (FR)"
"Y15-24","FR51",2009,19.4,"Pays de la Loire"
"Y15-24","FR52",2009,15.7,"Bretagne"
"Y15-24","FR53",2009,24.4,"Poitou-Charentes"
"Y15-24","FR6",2009,20.6,"Sud-Ouest (FR)"
"Y15-24","FR61",2009,21.9,"Aquitaine"
"Y15-24","FR62",2009,20.7,"Midi-Pyrénées"
"Y15-24","FR63",2009,NA,"Limousin"
"Y15-24","FR7",2009,21.1,"Centre-Est (FR)"
"Y15-24","FR71",2009,21.8,"Rhône-Alpes"
"Y15-24","FR72",2009,17,"Auvergne"
"Y15-24","FR8",2009,27.7,"Méditerranée"
"Y15-24","FR81",2009,33.7,"Languedoc-Roussillon"
"Y15-24","FR82",2009,25.2,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2009,NA,"Corse"
"Y15-24","FR9",2009,51.2,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2009,59.3,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2009,57.6,"Martinique (NUTS 2010)"
"Y15-24","FR93",2009,37.6,"Guyane (NUTS 2010)"
"Y15-24","FR94",2009,49.6,"Réunion (NUTS 2010)"
"Y15-24","HR",2009,25.2,"Croatia"
"Y15-24","HR0",2009,25.2,"Hrvatska"
"Y15-24","HR03",2009,22.9,"Jadranska Hrvatska"
"Y15-24","HR04",2009,26.2,"Kontinentalna Hrvatska"
"Y15-24","HU",2009,26.4,"Hungary"
"Y15-24","HU1",2009,18.6,"Közép-Magyarország"
"Y15-24","HU10",2009,18.6,"Közép-Magyarország"
"Y15-24","HU2",2009,25,"Dunántúl"
"Y15-24","HU21",2009,21.7,"Közép-Dunántúl"
"Y15-24","HU22",2009,23.6,"Nyugat-Dunántúl"
"Y15-24","HU23",2009,30.8,"Dél-Dunántúl"
"Y15-24","HU3",2009,32.2,"Alföld és Észak"
"Y15-24","HU31",2009,35.5,"Észak-Magyarország"
"Y15-24","HU32",2009,32.6,"Észak-Alföld"
"Y15-24","HU33",2009,28.1,"Dél-Alföld"
"Y15-24","IE",2009,24,"Ireland"
"Y15-24","IE0",2009,24,"Éire/Ireland"
"Y15-24","IE01",2009,27.2,"Border, Midland and Western"
"Y15-24","IE02",2009,22.9,"Southern and Eastern"
"Y15-24","IS",2009,15.9,"Iceland"
"Y15-24","IS0",2009,15.9,"Ísland"
"Y15-24","IS00",2009,15.9,"Ísland"
"Y15-24","IT",2009,25.3,"Italy"
"Y15-24","ITC",2009,20.1,"Nord-Ovest"
"Y15-24","ITC1",2009,24.3,"Piemonte"
"Y15-24","ITC2",2009,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2009,18.2,"Liguria"
"Y15-24","ITC4",2009,18.5,"Lombardia"
"Y15-24","ITF",2009,34,"Sud"
"Y15-24","ITF1",2009,24.4,"Abruzzo"
"Y15-24","ITF2",2009,27.1,"Molise"
"Y15-24","ITF3",2009,37.8,"Campania"
"Y15-24","ITF4",2009,32.7,"Puglia"
"Y15-24","ITF5",2009,38.3,"Basilicata"
"Y15-24","ITF6",2009,31.8,"Calabria"
"Y15-24","ITG",2009,39.7,"Isole"
"Y15-24","ITG1",2009,38.3,"Sicilia"
"Y15-24","ITG2",2009,44,"Sardegna"
"Y15-24","ITH",2009,15.3,"Nord-Est"
"Y15-24","ITH1",2009,8.9,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2009,11.6,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2009,14.3,"Veneto"
"Y15-24","ITH4",2009,18.2,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2009,17.8,"Emilia-Romagna"
"Y15-24","ITI",2009,24.4,"Centro (IT)"
"Y15-24","ITI1",2009,17.3,"Toscana"
"Y15-24","ITI2",2009,19,"Umbria"
"Y15-24","ITI3",2009,22.6,"Marche"
"Y15-24","ITI4",2009,30.4,"Lazio"
"Y15-24","LT",2009,29.6,"Lithuania"
"Y15-24","LT0",2009,29.6,"Lietuva"
"Y15-24","LT00",2009,29.6,"Lietuva"
"Y15-24","LU",2009,17.2,"Luxembourg"
"Y15-24","LU0",2009,17.2,"Luxembourg"
"Y15-24","LU00",2009,17.2,"Luxembourg"
"Y15-24","LV",2009,33.3,"Latvia"
"Y15-24","LV0",2009,33.3,"Latvija"
"Y15-24","LV00",2009,33.3,"Latvija"
"Y15-24","MK",2009,55.1,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2009,55.1,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2009,55.1,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2009,14.5,"Malta"
"Y15-24","MT0",2009,14.5,"Malta"
"Y15-24","MT00",2009,14.5,"Malta"
"Y15-24","NL",2009,6.6,"Netherlands"
"Y15-24","NL1",2009,8,"Noord-Nederland"
"Y15-24","NL11",2009,9.2,"Groningen"
"Y15-24","NL12",2009,7.3,"Friesland (NL)"
"Y15-24","NL13",2009,7.1,"Drenthe"
"Y15-24","NL2",2009,5.8,"Oost-Nederland"
"Y15-24","NL21",2009,5.6,"Overijssel"
"Y15-24","NL22",2009,5.4,"Gelderland"
"Y15-24","NL23",2009,8.3,"Flevoland"
"Y15-24","NL3",2009,6.6,"West-Nederland"
"Y15-24","NL31",2009,5.7,"Utrecht"
"Y15-24","NL32",2009,6.1,"Noord-Holland"
"Y15-24","NL33",2009,7.5,"Zuid-Holland"
"Y15-24","NL34",2009,NA,"Zeeland"
"Y15-24","NL4",2009,6.9,"Zuid-Nederland"
"Y15-24","NL41",2009,6.3,"Noord-Brabant"
"Y15-24","NL42",2009,8.4,"Limburg (NL)"
"Y15-24","NO",2009,9.2,"Norway"
"Y15-24","NO0",2009,9.2,"Norge"
"Y15-24","NO01",2009,10.8,"Oslo og Akershus"
"Y15-24","NO02",2009,8.4,"Hedmark og Oppland"
"Y15-24","NO03",2009,10.4,"Sør-Østlandet"
"Y15-24","NO04",2009,4.7,"Agder og Rogaland"
"Y15-24","NO05",2009,7.7,"Vestlandet"
"Y15-24","NO06",2009,10.4,"Trøndelag"
"Y15-24","NO07",2009,12.6,"Nord-Norge"
"Y15-24","PL",2009,20.6,"Poland"
"Y15-24","PL1",2009,16.2,"Region Centralny"
"Y15-24","PL11",2009,19.1,"Lódzkie"
"Y15-24","PL12",2009,14.9,"Mazowieckie"
"Y15-24","PL2",2009,20.9,"Region Poludniowy"
"Y15-24","PL21",2009,24.2,"Malopolskie"
"Y15-24","PL22",2009,18.3,"Slaskie"
"Y15-24","PL3",2009,26.4,"Region Wschodni"
"Y15-24","PL31",2009,26.9,"Lubelskie"
"Y15-24","PL32",2009,33.1,"Podkarpackie"
"Y15-24","PL33",2009,23.9,"Swietokrzyskie"
"Y15-24","PL34",2009,17.4,"Podlaskie"
"Y15-24","PL4",2009,20.1,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2009,17.8,"Wielkopolskie"
"Y15-24","PL42",2009,24.5,"Zachodniopomorskie"
"Y15-24","PL43",2009,23.5,"Lubuskie"
"Y15-24","PL5",2009,22.6,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2009,23.3,"Dolnoslaskie"
"Y15-24","PL52",2009,20.3,"Opolskie"
"Y15-24","PL6",2009,19.1,"Region Pólnocny"
"Y15-24","PL61",2009,21.5,"Kujawsko-Pomorskie"
"Y15-24","PL62",2009,18.8,"Warminsko-Mazurskie"
"Y15-24","PL63",2009,16.2,"Pomorskie"
"Y15-24","PT",2009,20.3,"Portugal"
"Y15-24","PT1",2009,20.5,"Continente"
"Y15-24","PT11",2009,22.2,"Norte"
"Y15-24","PT15",2009,24.8,"Algarve"
"Y15-24","PT16",2009,16.6,"Centro (PT)"
"Y15-24","PT17",2009,19,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2009,23.9,"Alentejo"
"Y15-24","PT2",2009,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2009,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2009,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2009,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2009,20.8,"Romania"
"Y15-24","RO1",2009,23.8,"Macroregiunea unu"
"Y15-24","RO11",2009,16.8,"Nord-Vest"
"Y15-24","RO12",2009,30.2,"Centru"
"Y15-24","RO2",2009,18.4,"Macroregiunea doi"
"Y15-24","RO21",2009,16.2,"Nord-Est"
"Y15-24","RO22",2009,21.8,"Sud-Est"
"Y15-24","RO3",2009,21.5,"Macroregiunea trei"
"Y15-24","RO31",2009,23.6,"Sud - Muntenia"
"Y15-24","RO32",2009,16.9,"Bucuresti - Ilfov"
"Y15-24","RO4",2009,20.1,"Macroregiunea patru"
"Y15-24","RO41",2009,20.3,"Sud-Vest Oltenia"
"Y15-24","RO42",2009,19.7,"Vest"
"Y15-24","SE",2009,25,"Sweden"
"Y15-24","SE1",2009,24,"Östra Sverige"
"Y15-24","SE11",2009,22.1,"Stockholm"
"Y15-24","SE12",2009,26.2,"Östra Mellansverige"
"Y15-24","SE2",2009,25.3,"Södra Sverige"
"Y15-24","SE21",2009,26.6,"Småland med öarna"
"Y15-24","SE22",2009,25.3,"Sydsverige"
"Y15-24","SE23",2009,24.8,"Västsverige"
"Y15-24","SE3",2009,26.4,"Norra Sverige"
"Y15-24","SE31",2009,25.8,"Norra Mellansverige"
"Y15-24","SE32",2009,30.8,"Mellersta Norrland"
"Y15-24","SE33",2009,24.5,"Övre Norrland"
"Y15-24","SI",2009,13.6,"Slovenia"
"Y15-24","SI0",2009,13.6,"Slovenija"
"Y15-24","SI01",2009,15.5,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2009,11.6,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2009,27.3,"Slovakia"
"Y15-24","SK0",2009,27.3,"Slovensko"
"Y15-24","SK01",2009,9.7,"Bratislavský kraj"
"Y15-24","SK02",2009,22.6,"Západné Slovensko"
"Y15-24","SK03",2009,32.5,"Stredné Slovensko"
"Y15-24","SK04",2009,34.4,"Východné Slovensko"
"Y15-24","TR",2009,22.8,"Turkey"
"Y15-24","TR1",2009,25.4,"Istanbul"
"Y15-24","TR10",2009,25.4,"Istanbul"
"Y15-24","TR2",2009,20.9,"Bati Marmara"
"Y15-24","TR21",2009,25.6,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2009,15,"Balikesir, Çanakkale"
"Y15-24","TR3",2009,24.9,"Ege"
"Y15-24","TR31",2009,30.4,"Izmir"
"Y15-24","TR32",2009,22.6,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2009,19.7,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2009,23.3,"Dogu Marmara"
"Y15-24","TR41",2009,22.5,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2009,24.3,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2009,21.6,"Bati Anadolu"
"Y15-24","TR51",2009,26.2,"Ankara"
"Y15-24","TR52",2009,15.4,"Konya, Karaman"
"Y15-24","TR6",2009,25.9,"Akdeniz"
"Y15-24","TR61",2009,19.6,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2009,31.6,"Adana, Mersin"
"Y15-24","TR63",2009,22.5,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2009,24.8,"Orta Anadolu"
"Y15-24","TR71",2009,27.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2009,22.5,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2009,13.3,"Bati Karadeniz"
"Y15-24","TR81",2009,19.4,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2009,17,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2009,10.4,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2009,12.8,"Dogu Karadeniz"
"Y15-24","TR90",2009,12.8,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2009,13.8,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2009,13.1,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2009,14.3,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2009,26.8,"Ortadogu Anadolu"
"Y15-24","TRB1",2009,30.7,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2009,23.4,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2009,21.6,"Güneydogu Anadolu"
"Y15-24","TRC1",2009,20.4,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2009,22,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2009,23.3,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2009,19.1,"United Kingdom"
"Y15-24","UKC",2009,22.9,"North East (UK)"
"Y15-24","UKC1",2009,21.7,"Tees Valley and Durham"
"Y15-24","UKC2",2009,23.7,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2009,21,"North West (UK)"
"Y15-24","UKD1",2009,20.3,"Cumbria"
"Y15-24","UKD3",2009,21.1,"Greater Manchester"
"Y15-24","UKD4",2009,17.7,"Lancashire"
"Y15-24","UKD6",2009,17.8,"Cheshire"
"Y15-24","UKD7",2009,26.6,"Merseyside"
"Y15-24","UKE",2009,20.2,"Yorkshire and The Humber"
"Y15-24","UKE1",2009,24.6,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2009,13.1,"North Yorkshire"
"Y15-24","UKE3",2009,22.3,"South Yorkshire"
"Y15-24","UKE4",2009,19.4,"West Yorkshire"
"Y15-24","UKF",2009,17.3,"East Midlands (UK)"
"Y15-24","UKF1",2009,15,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2009,18.2,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2009,21.7,"Lincolnshire"
"Y15-24","UKG",2009,24,"West Midlands (UK)"
"Y15-24","UKG1",2009,19.8,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2009,17.5,"Shropshire and Staffordshire"
"Y15-24","UKG3",2009,29.9,"West Midlands"
"Y15-24","UKH",2009,16.6,"East of England"
"Y15-24","UKH1",2009,17.3,"East Anglia"
"Y15-24","UKH2",2009,16.1,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2009,16,"Essex"
"Y15-24","UKI",2009,23,"London"
"Y15-24","UKI1",2009,25,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2009,21.6,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2009,16.2,"South East (UK)"
"Y15-24","UKJ1",2009,15.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2009,15.5,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2009,13.8,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2009,20.6,"Kent"
"Y15-24","UKK",2009,15.3,"South West (UK)"
"Y15-24","UKK1",2009,16.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2009,11.4,"Dorset and Somerset"
"Y15-24","UKK3",2009,12.2,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2009,18.4,"Devon"
"Y15-24","UKL",2009,19.9,"Wales"
"Y15-24","UKL1",2009,21.9,"West Wales and The Valleys"
"Y15-24","UKL2",2009,16,"East Wales"
"Y15-24","UKM",2009,16.6,"Scotland"
"Y15-24","UKM2",2009,20.5,"Eastern Scotland"
"Y15-24","UKM3",2009,15.9,"South Western Scotland"
"Y15-24","UKM5",2009,8.2,"North Eastern Scotland"
"Y15-24","UKM6",2009,NA,"Highlands and Islands"
"Y15-24","UKN",2009,16.7,"Northern Ireland (UK)"
"Y15-24","UKN0",2009,16.7,"Northern Ireland (UK)"
"Y20-64","AT",2009,5,"Austria"
"Y20-64","AT1",2009,6.2,"Ostösterreich"
"Y20-64","AT11",2009,4.8,"Burgenland (AT)"
"Y20-64","AT12",2009,4.3,"Niederösterreich"
"Y20-64","AT13",2009,8.3,"Wien"
"Y20-64","AT2",2009,4.6,"Südösterreich"
"Y20-64","AT21",2009,4.5,"Kärnten"
"Y20-64","AT22",2009,4.7,"Steiermark"
"Y20-64","AT3",2009,3.8,"Westösterreich"
"Y20-64","AT31",2009,4,"Oberösterreich"
"Y20-64","AT32",2009,3.2,"Salzburg"
"Y20-64","AT33",2009,3,"Tirol"
"Y20-64","AT34",2009,5.1,"Vorarlberg"
"Y20-64","BE",2009,7.7,"Belgium"
"Y20-64","BE1",2009,15.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2009,15.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2009,4.7,"Vlaams Gewest"
"Y20-64","BE21",2009,5.6,"Prov. Antwerpen"
"Y20-64","BE22",2009,5.1,"Prov. Limburg (BE)"
"Y20-64","BE23",2009,4.1,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2009,4.7,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2009,4.1,"Prov. West-Vlaanderen"
"Y20-64","BE3",2009,10.9,"Région wallonne"
"Y20-64","BE31",2009,6.6,"Prov. Brabant Wallon"
"Y20-64","BE32",2009,12.7,"Prov. Hainaut"
"Y20-64","BE33",2009,11.9,"Prov. Liège"
"Y20-64","BE34",2009,7.2,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2009,9.2,"Prov. Namur"
"Y20-64","BG",2009,6.6,"Bulgaria"
"Y20-64","BG3",2009,8.1,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2009,7.9,"Severozapaden"
"Y20-64","BG32",2009,7.9,"Severen tsentralen"
"Y20-64","BG33",2009,10.1,"Severoiztochen"
"Y20-64","BG34",2009,6.4,"Yugoiztochen"
"Y20-64","BG4",2009,5.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2009,4,"Yugozapaden"
"Y20-64","BG42",2009,6.9,"Yuzhen tsentralen"
"Y20-64","CH",2009,4,"Switzerland"
"Y20-64","CH0",2009,4,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2009,5.4,"Région lémanique"
"Y20-64","CH02",2009,3.5,"Espace Mittelland"
"Y20-64","CH03",2009,4.5,"Nordwestschweiz"
"Y20-64","CH04",2009,3.7,"Zürich"
"Y20-64","CH05",2009,3.4,"Ostschweiz"
"Y20-64","CH06",2009,2.6,"Zentralschweiz"
"Y20-64","CH07",2009,5,"Ticino"
"Y20-64","CY",2009,5.4,"Cyprus"
"Y20-64","CY0",2009,5.4,"Kypros"
"Y20-64","CY00",2009,5.4,"Kypros"
"Y20-64","CZ",2009,6.5,"Czech Republic"
"Y20-64","CZ0",2009,6.5,"Ceská republika"
"Y20-64","CZ01",2009,3,"Praha"
"Y20-64","CZ02",2009,4.1,"Strední Cechy"
"Y20-64","CZ03",2009,5,"Jihozápad"
"Y20-64","CZ04",2009,9.8,"Severozápad"
"Y20-64","CZ05",2009,7.1,"Severovýchod"
"Y20-64","CZ06",2009,6.4,"Jihovýchod"
"Y20-64","CZ07",2009,7.3,"Strední Morava"
"Y20-64","CZ08",2009,9.5,"Moravskoslezsko"
"Y20-64","DE",2009,7.7,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2009,5.1,"Baden-Württemberg"
"Y20-64","DE11",2009,5.1,"Stuttgart"
"Y20-64","DE12",2009,5.5,"Karlsruhe"
"Y20-64","DE13",2009,4.3,"Freiburg"
"Y20-64","DE14",2009,5.1,"Tübingen"
"Y20-64","DE2",2009,5,"Bayern"
"Y20-64","DE21",2009,4.2,"Oberbayern"
"Y20-64","DE22",2009,5,"Niederbayern"
"Y20-64","DE23",2009,4.9,"Oberpfalz"
"Y20-64","DE24",2009,6.6,"Oberfranken"
"Y20-64","DE25",2009,6.4,"Mittelfranken"
"Y20-64","DE26",2009,5.5,"Unterfranken"
"Y20-64","DE27",2009,4.6,"Schwaben"
"Y20-64","DE3",2009,13.8,"Berlin"
"Y20-64","DE30",2009,13.8,"Berlin"
"Y20-64","DE4",2009,11.3,"Brandenburg"
"Y20-64","DE40",2009,11.3,"Brandenburg"
"Y20-64","DE5",2009,9.1,"Bremen"
"Y20-64","DE50",2009,9.1,"Bremen"
"Y20-64","DE6",2009,7.2,"Hamburg"
"Y20-64","DE60",2009,7.2,"Hamburg"
"Y20-64","DE7",2009,6.3,"Hessen"
"Y20-64","DE71",2009,6.1,"Darmstadt"
"Y20-64","DE72",2009,6.6,"Gießen"
"Y20-64","DE73",2009,6.5,"Kassel"
"Y20-64","DE8",2009,14.1,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2009,14.1,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2009,6.9,"Niedersachsen"
"Y20-64","DE91",2009,8.5,"Braunschweig"
"Y20-64","DE92",2009,8,"Hannover"
"Y20-64","DE93",2009,5.4,"Lüneburg"
"Y20-64","DE94",2009,5.9,"Weser-Ems"
"Y20-64","DEA",2009,7.8,"Nordrhein-Westfalen"
"Y20-64","DEA1",2009,7.6,"Düsseldorf"
"Y20-64","DEA2",2009,7.1,"Köln"
"Y20-64","DEA3",2009,7.3,"Münster"
"Y20-64","DEA4",2009,7.7,"Detmold"
"Y20-64","DEA5",2009,9.2,"Arnsberg"
"Y20-64","DEB",2009,5.8,"Rheinland-Pfalz"
"Y20-64","DEB1",2009,6.6,"Koblenz"
"Y20-64","DEB2",2009,4.5,"Trier"
"Y20-64","DEB3",2009,5.5,"Rheinhessen-Pfalz"
"Y20-64","DEC",2009,8.3,"Saarland"
"Y20-64","DEC0",2009,8.3,"Saarland"
"Y20-64","DED",2009,12.6,"Sachsen"
"Y20-64","DED2",2009,12,"Dresden"
"Y20-64","DED4",2009,12.8,"Chemnitz"
"Y20-64","DED5",2009,13.1,"Leipzig"
"Y20-64","DEE",2009,13.7,"Sachsen-Anhalt"
"Y20-64","DEE0",2009,13.7,"Sachsen-Anhalt"
"Y20-64","DEF",2009,7.4,"Schleswig-Holstein"
"Y20-64","DEF0",2009,7.4,"Schleswig-Holstein"
"Y20-64","DEG",2009,10.8,"Thüringen"
"Y20-64","DEG0",2009,10.8,"Thüringen"
"Y20-64","DK",2009,5.5,"Denmark"
"Y20-64","DK0",2009,5.5,"Danmark"
"Y20-64","DK01",2009,5.6,"Hovedstaden"
"Y20-64","DK02",2009,4.7,"Sjælland"
"Y20-64","DK03",2009,5.5,"Syddanmark"
"Y20-64","DK04",2009,5.4,"Midtjylland"
"Y20-64","DK05",2009,6.5,"Nordjylland"
"Y20-64","EA17",2009,9.2,"Euro area (17 countries)"
"Y20-64","EA18",2009,9.3,"Euro area (18 countries)"
"Y20-64","EA19",2009,9.3,"Euro area (19 countries)"
"Y20-64","EE",2009,13.3,"Estonia"
"Y20-64","EE0",2009,13.3,"Eesti"
"Y20-64","EE00",2009,13.3,"Eesti"
"Y20-64","EL",2009,9.5,"Greece"
"Y20-64","EL1",2009,10.3,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2009,11,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2009,10,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2009,12.5,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2009,9.5,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2009,9.6,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2009,11.3,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2009,9.3,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2009,9.7,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2009,10.4,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2009,8,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2009,8.9,"Attiki"
"Y20-64","EL30",2009,8.9,"Attiki"
"Y20-64","EL4",2009,9.5,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2009,6.4,"Voreio Aigaio"
"Y20-64","EL42",2009,12,"Notio Aigaio"
"Y20-64","EL43",2009,9,"Kriti"
"Y20-64","ES",2009,17.2,"Spain"
"Y20-64","ES1",2009,12.3,"Noroeste (ES)"
"Y20-64","ES11",2009,12.1,"Galicia"
"Y20-64","ES12",2009,13,"Principado de Asturias"
"Y20-64","ES13",2009,11.7,"Cantabria"
"Y20-64","ES2",2009,11.5,"Noreste (ES)"
"Y20-64","ES21",2009,11.1,"País Vasco"
"Y20-64","ES22",2009,10.1,"Comunidad Foral de Navarra"
"Y20-64","ES23",2009,11.8,"La Rioja"
"Y20-64","ES24",2009,12.6,"Aragón"
"Y20-64","ES3",2009,13.3,"Comunidad de Madrid"
"Y20-64","ES30",2009,13.3,"Comunidad de Madrid"
"Y20-64","ES4",2009,16.3,"Centro (ES)"
"Y20-64","ES41",2009,13.5,"Castilla y León"
"Y20-64","ES42",2009,18,"Castilla-la Mancha"
"Y20-64","ES43",2009,19.8,"Extremadura"
"Y20-64","ES5",2009,17.3,"Este (ES)"
"Y20-64","ES51",2009,15.5,"Cataluña"
"Y20-64","ES52",2009,20,"Comunidad Valenciana"
"Y20-64","ES53",2009,17.3,"Illes Balears"
"Y20-64","ES6",2009,23.6,"Sur (ES)"
"Y20-64","ES61",2009,24.4,"Andalucía"
"Y20-64","ES62",2009,19.5,"Región de Murcia"
"Y20-64","ES63",2009,18.1,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2009,23.6,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2009,25.5,"Canarias (ES)"
"Y20-64","ES70",2009,25.5,"Canarias (ES)"
"Y20-64","EU15",2009,8.7,"European Union (15 countries)"
"Y20-64","EU27",2009,8.6,"European Union (27 countries)"
"Y20-64","EU28",2009,8.6,"European Union (28 countries)"
"Y20-64","FI",2009,7.4,"Finland"
"Y20-64","FI1",2009,7.5,"Manner-Suomi"
"Y20-64","FI19",2009,8.3,"Länsi-Suomi"
"Y20-64","FI1B",2009,5.4,"Helsinki-Uusimaa"
"Y20-64","FI1C",2009,7.3,"Etelä-Suomi"
"Y20-64","FI1D",2009,9.6,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2009,NA,"Åland"
"Y20-64","FI20",2009,NA,"Åland"
"Y20-64","FR",2009,8.7,"France"
"Y20-64","FR1",2009,7.8,"Île de France"
"Y20-64","FR10",2009,7.8,"Île de France"
"Y20-64","FR2",2009,7.9,"Bassin Parisien"
"Y20-64","FR21",2009,8.8,"Champagne-Ardenne"
"Y20-64","FR22",2009,9.9,"Picardie"
"Y20-64","FR23",2009,9.3,"Haute-Normandie"
"Y20-64","FR24",2009,6.2,"Centre (FR)"
"Y20-64","FR25",2009,6.5,"Basse-Normandie"
"Y20-64","FR26",2009,7.1,"Bourgogne"
"Y20-64","FR3",2009,12.4,"Nord - Pas-de-Calais"
"Y20-64","FR30",2009,12.4,"Nord - Pas-de-Calais"
"Y20-64","FR4",2009,9,"Est (FR)"
"Y20-64","FR41",2009,10.3,"Lorraine"
"Y20-64","FR42",2009,7.8,"Alsace"
"Y20-64","FR43",2009,8.3,"Franche-Comté"
"Y20-64","FR5",2009,6.7,"Ouest (FR)"
"Y20-64","FR51",2009,7.2,"Pays de la Loire"
"Y20-64","FR52",2009,5.3,"Bretagne"
"Y20-64","FR53",2009,8,"Poitou-Charentes"
"Y20-64","FR6",2009,7.9,"Sud-Ouest (FR)"
"Y20-64","FR61",2009,8,"Aquitaine"
"Y20-64","FR62",2009,8.3,"Midi-Pyrénées"
"Y20-64","FR63",2009,6,"Limousin"
"Y20-64","FR7",2009,7.7,"Centre-Est (FR)"
"Y20-64","FR71",2009,7.8,"Rhône-Alpes"
"Y20-64","FR72",2009,7.1,"Auvergne"
"Y20-64","FR8",2009,9.9,"Méditerranée"
"Y20-64","FR81",2009,12.5,"Languedoc-Roussillon"
"Y20-64","FR82",2009,8.7,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2009,NA,"Corse"
"Y20-64","FR9",2009,23.7,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2009,22.9,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2009,21.2,"Martinique (NUTS 2010)"
"Y20-64","FR93",2009,19.7,"Guyane (NUTS 2010)"
"Y20-64","FR94",2009,26.2,"Réunion (NUTS 2010)"
"Y20-64","HR",2009,8.8,"Croatia"
"Y20-64","HR0",2009,8.8,"Hrvatska"
"Y20-64","HR03",2009,9.2,"Jadranska Hrvatska"
"Y20-64","HR04",2009,8.7,"Kontinentalna Hrvatska"
"Y20-64","HU",2009,9.9,"Hungary"
"Y20-64","HU1",2009,6.4,"Közép-Magyarország"
"Y20-64","HU10",2009,6.4,"Közép-Magyarország"
"Y20-64","HU2",2009,9.4,"Dunántúl"
"Y20-64","HU21",2009,9,"Közép-Dunántúl"
"Y20-64","HU22",2009,8.6,"Nyugat-Dunántúl"
"Y20-64","HU23",2009,10.9,"Dél-Dunántúl"
"Y20-64","HU3",2009,13.1,"Alföld és Észak"
"Y20-64","HU31",2009,15,"Észak-Magyarország"
"Y20-64","HU32",2009,13.9,"Észak-Alföld"
"Y20-64","HU33",2009,10.5,"Dél-Alföld"
"Y20-64","IE",2009,11.7,"Ireland"
"Y20-64","IE0",2009,11.7,"Éire/Ireland"
"Y20-64","IE01",2009,13,"Border, Midland and Western"
"Y20-64","IE02",2009,11.2,"Southern and Eastern"
"Y20-64","IS",2009,6.6,"Iceland"
"Y20-64","IS0",2009,6.6,"Ísland"
"Y20-64","IS00",2009,6.6,"Ísland"
"Y20-64","IT",2009,7.5,"Italy"
"Y20-64","ITC",2009,5.5,"Nord-Ovest"
"Y20-64","ITC1",2009,6.5,"Piemonte"
"Y20-64","ITC2",2009,4.3,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2009,5.8,"Liguria"
"Y20-64","ITC4",2009,5,"Lombardia"
"Y20-64","ITF",2009,11.5,"Sud"
"Y20-64","ITF1",2009,7.7,"Abruzzo"
"Y20-64","ITF2",2009,8.8,"Molise"
"Y20-64","ITF3",2009,12.5,"Campania"
"Y20-64","ITF4",2009,12.2,"Puglia"
"Y20-64","ITF5",2009,10.9,"Basilicata"
"Y20-64","ITF6",2009,11.1,"Calabria"
"Y20-64","ITG",2009,13.1,"Isole"
"Y20-64","ITG1",2009,13.2,"Sicilia"
"Y20-64","ITG2",2009,12.9,"Sardegna"
"Y20-64","ITH",2009,4.4,"Nord-Est"
"Y20-64","ITH1",2009,2.7,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2009,3.3,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2009,4.4,"Veneto"
"Y20-64","ITH4",2009,5,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2009,4.6,"Emilia-Romagna"
"Y20-64","ITI",2009,7,"Centro (IT)"
"Y20-64","ITI1",2009,5.6,"Toscana"
"Y20-64","ITI2",2009,6.4,"Umbria"
"Y20-64","ITI3",2009,6.4,"Marche"
"Y20-64","ITI4",2009,8.2,"Lazio"
"Y20-64","LT",2009,13.7,"Lithuania"
"Y20-64","LT0",2009,13.7,"Lietuva"
"Y20-64","LT00",2009,13.7,"Lietuva"
"Y20-64","LU",2009,4.9,"Luxembourg"
"Y20-64","LU0",2009,4.9,"Luxembourg"
"Y20-64","LU00",2009,4.9,"Luxembourg"
"Y20-64","LV",2009,17.3,"Latvia"
"Y20-64","LV0",2009,17.3,"Latvija"
"Y20-64","LV00",2009,17.3,"Latvija"
"Y20-64","MK",2009,31.7,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2009,31.7,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2009,31.7,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2009,5.9,"Malta"
"Y20-64","MT0",2009,5.9,"Malta"
"Y20-64","MT00",2009,5.9,"Malta"
"Y20-64","NL",2009,3,"Netherlands"
"Y20-64","NL1",2009,3.7,"Noord-Nederland"
"Y20-64","NL11",2009,4.3,"Groningen"
"Y20-64","NL12",2009,3.1,"Friesland (NL)"
"Y20-64","NL13",2009,3.9,"Drenthe"
"Y20-64","NL2",2009,2.8,"Oost-Nederland"
"Y20-64","NL21",2009,3.3,"Overijssel"
"Y20-64","NL22",2009,2.4,"Gelderland"
"Y20-64","NL23",2009,2.9,"Flevoland"
"Y20-64","NL3",2009,2.9,"West-Nederland"
"Y20-64","NL31",2009,2.6,"Utrecht"
"Y20-64","NL32",2009,2.9,"Noord-Holland"
"Y20-64","NL33",2009,3.1,"Zuid-Holland"
"Y20-64","NL34",2009,2,"Zeeland"
"Y20-64","NL4",2009,3.2,"Zuid-Nederland"
"Y20-64","NL41",2009,2.9,"Noord-Brabant"
"Y20-64","NL42",2009,4,"Limburg (NL)"
"Y20-64","NO",2009,2.6,"Norway"
"Y20-64","NO0",2009,2.6,"Norge"
"Y20-64","NO01",2009,3.2,"Oslo og Akershus"
"Y20-64","NO02",2009,2,"Hedmark og Oppland"
"Y20-64","NO03",2009,2.9,"Sør-Østlandet"
"Y20-64","NO04",2009,2.1,"Agder og Rogaland"
"Y20-64","NO05",2009,2,"Vestlandet"
"Y20-64","NO06",2009,3.1,"Trøndelag"
"Y20-64","NO07",2009,2.8,"Nord-Norge"
"Y20-64","PL",2009,8.1,"Poland"
"Y20-64","PL1",2009,6.4,"Region Centralny"
"Y20-64","PL11",2009,7.5,"Lódzkie"
"Y20-64","PL12",2009,5.8,"Mazowieckie"
"Y20-64","PL2",2009,7.1,"Region Poludniowy"
"Y20-64","PL21",2009,7.8,"Malopolskie"
"Y20-64","PL22",2009,6.6,"Slaskie"
"Y20-64","PL3",2009,9.7,"Region Wschodni"
"Y20-64","PL31",2009,9.8,"Lubelskie"
"Y20-64","PL32",2009,10.1,"Podkarpackie"
"Y20-64","PL33",2009,11,"Swietokrzyskie"
"Y20-64","PL34",2009,7,"Podlaskie"
"Y20-64","PL4",2009,8.4,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2009,7.2,"Wielkopolskie"
"Y20-64","PL42",2009,10,"Zachodniopomorskie"
"Y20-64","PL43",2009,9.3,"Lubuskie"
"Y20-64","PL5",2009,9.9,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2009,9.9,"Dolnoslaskie"
"Y20-64","PL52",2009,9.8,"Opolskie"
"Y20-64","PL6",2009,8.4,"Region Pólnocny"
"Y20-64","PL61",2009,10.2,"Kujawsko-Pomorskie"
"Y20-64","PL62",2009,8.4,"Warminsko-Mazurskie"
"Y20-64","PL63",2009,6.4,"Pomorskie"
"Y20-64","PT",2009,9.7,"Portugal"
"Y20-64","PT1",2009,9.9,"Continente"
"Y20-64","PT11",2009,11.2,"Norte"
"Y20-64","PT15",2009,10.3,"Algarve"
"Y20-64","PT16",2009,7.5,"Centro (PT)"
"Y20-64","PT17",2009,9.8,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2009,10.7,"Alentejo"
"Y20-64","PT2",2009,6.5,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2009,6.5,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2009,7.6,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2009,7.6,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2009,6.7,"Romania"
"Y20-64","RO1",2009,7.7,"Macroregiunea unu"
"Y20-64","RO11",2009,5.5,"Nord-Vest"
"Y20-64","RO12",2009,10,"Centru"
"Y20-64","RO2",2009,6.5,"Macroregiunea doi"
"Y20-64","RO21",2009,6.1,"Nord-Est"
"Y20-64","RO22",2009,7.2,"Sud-Est"
"Y20-64","RO3",2009,6.1,"Macroregiunea trei"
"Y20-64","RO31",2009,7.9,"Sud - Muntenia"
"Y20-64","RO32",2009,3.6,"Bucuresti - Ilfov"
"Y20-64","RO4",2009,6.4,"Macroregiunea patru"
"Y20-64","RO41",2009,7.1,"Sud-Vest Oltenia"
"Y20-64","RO42",2009,5.7,"Vest"
"Y20-64","SE",2009,7.3,"Sweden"
"Y20-64","SE1",2009,6.8,"Östra Sverige"
"Y20-64","SE11",2009,5.7,"Stockholm"
"Y20-64","SE12",2009,8.3,"Östra Mellansverige"
"Y20-64","SE2",2009,7.4,"Södra Sverige"
"Y20-64","SE21",2009,7,"Småland med öarna"
"Y20-64","SE22",2009,7.7,"Sydsverige"
"Y20-64","SE23",2009,7.4,"Västsverige"
"Y20-64","SE3",2009,8,"Norra Sverige"
"Y20-64","SE31",2009,8.4,"Norra Mellansverige"
"Y20-64","SE32",2009,7.4,"Mellersta Norrland"
"Y20-64","SE33",2009,7.9,"Övre Norrland"
"Y20-64","SI",2009,5.8,"Slovenia"
"Y20-64","SI0",2009,5.8,"Slovenija"
"Y20-64","SI01",2009,6.8,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2009,4.8,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2009,11.7,"Slovakia"
"Y20-64","SK0",2009,11.7,"Slovensko"
"Y20-64","SK01",2009,4.6,"Bratislavský kraj"
"Y20-64","SK02",2009,9.7,"Západné Slovensko"
"Y20-64","SK03",2009,14.1,"Stredné Slovensko"
"Y20-64","SK04",2009,15.3,"Východné Slovensko"
"Y20-64","TR",2009,12.2,"Turkey"
"Y20-64","TR1",2009,15.2,"Istanbul"
"Y20-64","TR10",2009,15.2,"Istanbul"
"Y20-64","TR2",2009,9.1,"Bati Marmara"
"Y20-64","TR21",2009,11.2,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2009,7,"Balikesir, Çanakkale"
"Y20-64","TR3",2009,12.6,"Ege"
"Y20-64","TR31",2009,14.8,"Izmir"
"Y20-64","TR32",2009,12.7,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2009,9.1,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2009,12.4,"Dogu Marmara"
"Y20-64","TR41",2009,12.3,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2009,12.5,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2009,10.6,"Bati Anadolu"
"Y20-64","TR51",2009,11.6,"Ankara"
"Y20-64","TR52",2009,8.6,"Konya, Karaman"
"Y20-64","TR6",2009,15.1,"Akdeniz"
"Y20-64","TR61",2009,10,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2009,19.3,"Adana, Mersin"
"Y20-64","TR63",2009,15,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2009,12.2,"Orta Anadolu"
"Y20-64","TR71",2009,13.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2009,11,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2009,6.6,"Bati Karadeniz"
"Y20-64","TR81",2009,6.7,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2009,8.6,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2009,6.1,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2009,4.3,"Dogu Karadeniz"
"Y20-64","TR90",2009,4.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2009,6.6,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2009,6.3,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2009,6.9,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2009,14,"Ortadogu Anadolu"
"Y20-64","TRB1",2009,14.3,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2009,13.6,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2009,14.7,"Güneydogu Anadolu"
"Y20-64","TRC1",2009,14.1,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2009,16.1,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2009,13.2,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2009,6.6,"United Kingdom"
"Y20-64","UKC",2009,7.7,"North East (UK)"
"Y20-64","UKC1",2009,6.9,"Tees Valley and Durham"
"Y20-64","UKC2",2009,8.4,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2009,7.3,"North West (UK)"
"Y20-64","UKD1",2009,5.1,"Cumbria"
"Y20-64","UKD3",2009,8.4,"Greater Manchester"
"Y20-64","UKD4",2009,6.4,"Lancashire"
"Y20-64","UKD6",2009,4.8,"Cheshire"
"Y20-64","UKD7",2009,8.4,"Merseyside"
"Y20-64","UKE",2009,7.4,"Yorkshire and The Humber"
"Y20-64","UKE1",2009,7.9,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2009,4.7,"North Yorkshire"
"Y20-64","UKE3",2009,8.5,"South Yorkshire"
"Y20-64","UKE4",2009,7.5,"West Yorkshire"
"Y20-64","UKF",2009,6.2,"East Midlands (UK)"
"Y20-64","UKF1",2009,6.3,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2009,6.4,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2009,5.1,"Lincolnshire"
"Y20-64","UKG",2009,8.6,"West Midlands (UK)"
"Y20-64","UKG1",2009,5.4,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2009,6.4,"Shropshire and Staffordshire"
"Y20-64","UKG3",2009,11.7,"West Midlands"
"Y20-64","UKH",2009,5.2,"East of England"
"Y20-64","UKH1",2009,4.6,"East Anglia"
"Y20-64","UKH2",2009,5.4,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2009,5.9,"Essex"
"Y20-64","UKI",2009,8,"London"
"Y20-64","UKI1",2009,8.6,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2009,7.6,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2009,5,"South East (UK)"
"Y20-64","UKJ1",2009,4.7,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2009,4.9,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2009,4.5,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2009,6.1,"Kent"
"Y20-64","UKK",2009,5.3,"South West (UK)"
"Y20-64","UKK1",2009,4.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2009,5.9,"Dorset and Somerset"
"Y20-64","UKK3",2009,4.5,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2009,6.2,"Devon"
"Y20-64","UKL",2009,7,"Wales"
"Y20-64","UKL1",2009,7.7,"West Wales and The Valleys"
"Y20-64","UKL2",2009,6,"East Wales"
"Y20-64","UKM",2009,5.9,"Scotland"
"Y20-64","UKM2",2009,6.3,"Eastern Scotland"
"Y20-64","UKM3",2009,6.7,"South Western Scotland"
"Y20-64","UKM5",2009,3.4,"North Eastern Scotland"
"Y20-64","UKM6",2009,3.4,"Highlands and Islands"
"Y20-64","UKN",2009,5.9,"Northern Ireland (UK)"
"Y20-64","UKN0",2009,5.9,"Northern Ireland (UK)"
"Y_GE15","AT",2009,5.3,"Austria"
"Y_GE15","AT1",2009,6.6,"Ostösterreich"
"Y_GE15","AT11",2009,5,"Burgenland (AT)"
"Y_GE15","AT12",2009,4.7,"Niederösterreich"
"Y_GE15","AT13",2009,8.7,"Wien"
"Y_GE15","AT2",2009,4.9,"Südösterreich"
"Y_GE15","AT21",2009,4.6,"Kärnten"
"Y_GE15","AT22",2009,5,"Steiermark"
"Y_GE15","AT3",2009,4.1,"Westösterreich"
"Y_GE15","AT31",2009,4.2,"Oberösterreich"
"Y_GE15","AT32",2009,3.6,"Salzburg"
"Y_GE15","AT33",2009,3.3,"Tirol"
"Y_GE15","AT34",2009,5.6,"Vorarlberg"
"Y_GE15","BE",2009,7.9,"Belgium"
"Y_GE15","BE1",2009,15.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2009,15.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2009,4.9,"Vlaams Gewest"
"Y_GE15","BE21",2009,5.7,"Prov. Antwerpen"
"Y_GE15","BE22",2009,5.4,"Prov. Limburg (BE)"
"Y_GE15","BE23",2009,4.2,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2009,4.9,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2009,4.3,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2009,11.2,"Région wallonne"
"Y_GE15","BE31",2009,6.9,"Prov. Brabant Wallon"
"Y_GE15","BE32",2009,13.2,"Prov. Hainaut"
"Y_GE15","BE33",2009,12.1,"Prov. Liège"
"Y_GE15","BE34",2009,7.4,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2009,9.4,"Prov. Namur"
"Y_GE15","BG",2009,6.8,"Bulgaria"
"Y_GE15","BG3",2009,8.3,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2009,8,"Severozapaden"
"Y_GE15","BG32",2009,8.4,"Severen tsentralen"
"Y_GE15","BG33",2009,10.4,"Severoiztochen"
"Y_GE15","BG34",2009,6.6,"Yugoiztochen"
"Y_GE15","BG4",2009,5.3,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2009,4.1,"Yugozapaden"
"Y_GE15","BG42",2009,7.3,"Yuzhen tsentralen"
"Y_GE15","CH",2009,4.1,"Switzerland"
"Y_GE15","CH0",2009,4.1,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2009,5.9,"Région lémanique"
"Y_GE15","CH02",2009,3.6,"Espace Mittelland"
"Y_GE15","CH03",2009,4.5,"Nordwestschweiz"
"Y_GE15","CH04",2009,3.8,"Zürich"
"Y_GE15","CH05",2009,3.4,"Ostschweiz"
"Y_GE15","CH06",2009,2.7,"Zentralschweiz"
"Y_GE15","CH07",2009,5.1,"Ticino"
"Y_GE15","CY",2009,5.4,"Cyprus"
"Y_GE15","CY0",2009,5.4,"Kypros"
"Y_GE15","CY00",2009,5.4,"Kypros"
"Y_GE15","CZ",2009,6.7,"Czech Republic"
"Y_GE15","CZ0",2009,6.7,"Ceská republika"
"Y_GE15","CZ01",2009,3.1,"Praha"
"Y_GE15","CZ02",2009,4.4,"Strední Cechy"
"Y_GE15","CZ03",2009,5.2,"Jihozápad"
"Y_GE15","CZ04",2009,10.3,"Severozápad"
"Y_GE15","CZ05",2009,7.3,"Severovýchod"
"Y_GE15","CZ06",2009,6.5,"Jihovýchod"
"Y_GE15","CZ07",2009,7.5,"Strední Morava"
"Y_GE15","CZ08",2009,9.7,"Moravskoslezsko"
"Y_GE15","DE",2009,7.7,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2009,5.1,"Baden-Württemberg"
"Y_GE15","DE11",2009,5.3,"Stuttgart"
"Y_GE15","DE12",2009,5.6,"Karlsruhe"
"Y_GE15","DE13",2009,4.4,"Freiburg"
"Y_GE15","DE14",2009,5,"Tübingen"
"Y_GE15","DE2",2009,5.1,"Bayern"
"Y_GE15","DE21",2009,4.2,"Oberbayern"
"Y_GE15","DE22",2009,5,"Niederbayern"
"Y_GE15","DE23",2009,5,"Oberpfalz"
"Y_GE15","DE24",2009,6.7,"Oberfranken"
"Y_GE15","DE25",2009,6.4,"Mittelfranken"
"Y_GE15","DE26",2009,5.7,"Unterfranken"
"Y_GE15","DE27",2009,4.7,"Schwaben"
"Y_GE15","DE3",2009,13.7,"Berlin"
"Y_GE15","DE30",2009,13.7,"Berlin"
"Y_GE15","DE4",2009,11.3,"Brandenburg"
"Y_GE15","DE40",2009,11.3,"Brandenburg"
"Y_GE15","DE5",2009,9.1,"Bremen"
"Y_GE15","DE50",2009,9.1,"Bremen"
"Y_GE15","DE6",2009,7.2,"Hamburg"
"Y_GE15","DE60",2009,7.2,"Hamburg"
"Y_GE15","DE7",2009,6.4,"Hessen"
"Y_GE15","DE71",2009,6.3,"Darmstadt"
"Y_GE15","DE72",2009,6.7,"Gießen"
"Y_GE15","DE73",2009,6.6,"Kassel"
"Y_GE15","DE8",2009,13.9,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2009,13.9,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2009,6.9,"Niedersachsen"
"Y_GE15","DE91",2009,8.5,"Braunschweig"
"Y_GE15","DE92",2009,7.9,"Hannover"
"Y_GE15","DE93",2009,5.4,"Lüneburg"
"Y_GE15","DE94",2009,5.9,"Weser-Ems"
"Y_GE15","DEA",2009,7.8,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2009,7.7,"Düsseldorf"
"Y_GE15","DEA2",2009,7.1,"Köln"
"Y_GE15","DEA3",2009,7.3,"Münster"
"Y_GE15","DEA4",2009,7.7,"Detmold"
"Y_GE15","DEA5",2009,9.2,"Arnsberg"
"Y_GE15","DEB",2009,6,"Rheinland-Pfalz"
"Y_GE15","DEB1",2009,6.7,"Koblenz"
"Y_GE15","DEB2",2009,4.6,"Trier"
"Y_GE15","DEB3",2009,5.8,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2009,8.4,"Saarland"
"Y_GE15","DEC0",2009,8.4,"Saarland"
"Y_GE15","DED",2009,12.5,"Sachsen"
"Y_GE15","DED2",2009,12,"Dresden"
"Y_GE15","DED4",2009,12.5,"Chemnitz"
"Y_GE15","DED5",2009,13.1,"Leipzig"
"Y_GE15","DEE",2009,13.7,"Sachsen-Anhalt"
"Y_GE15","DEE0",2009,13.7,"Sachsen-Anhalt"
"Y_GE15","DEF",2009,7.3,"Schleswig-Holstein"
"Y_GE15","DEF0",2009,7.3,"Schleswig-Holstein"
"Y_GE15","DEG",2009,10.7,"Thüringen"
"Y_GE15","DEG0",2009,10.7,"Thüringen"
"Y_GE15","DK",2009,6,"Denmark"
"Y_GE15","DK0",2009,6,"Danmark"
"Y_GE15","DK01",2009,6.2,"Hovedstaden"
"Y_GE15","DK02",2009,5.3,"Sjælland"
"Y_GE15","DK03",2009,6,"Syddanmark"
"Y_GE15","DK04",2009,5.8,"Midtjylland"
"Y_GE15","DK05",2009,6.9,"Nordjylland"
"Y_GE15","EA17",2009,9.5,"Euro area (17 countries)"
"Y_GE15","EA18",2009,9.5,"Euro area (18 countries)"
"Y_GE15","EA19",2009,9.6,"Euro area (19 countries)"
"Y_GE15","EE",2009,13.5,"Estonia"
"Y_GE15","EE0",2009,13.5,"Eesti"
"Y_GE15","EE00",2009,13.5,"Eesti"
"Y_GE15","EL",2009,9.6,"Greece"
"Y_GE15","EL1",2009,10.3,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2009,11.1,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2009,10.1,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2009,12.4,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2009,9.2,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2009,9.6,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2009,11.2,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2009,9.5,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2009,9.7,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2009,10.5,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2009,7.9,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2009,9.1,"Attiki"
"Y_GE15","EL30",2009,9.1,"Attiki"
"Y_GE15","EL4",2009,9.6,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2009,6.6,"Voreio Aigaio"
"Y_GE15","EL42",2009,12.3,"Notio Aigaio"
"Y_GE15","EL43",2009,9,"Kriti"
"Y_GE15","ES",2009,17.9,"Spain"
"Y_GE15","ES1",2009,12.6,"Noroeste (ES)"
"Y_GE15","ES11",2009,12.4,"Galicia"
"Y_GE15","ES12",2009,13.4,"Principado de Asturias"
"Y_GE15","ES13",2009,12,"Cantabria"
"Y_GE15","ES2",2009,11.9,"Noreste (ES)"
"Y_GE15","ES21",2009,11.3,"País Vasco"
"Y_GE15","ES22",2009,10.8,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2009,12.6,"La Rioja"
"Y_GE15","ES24",2009,13.1,"Aragón"
"Y_GE15","ES3",2009,13.9,"Comunidad de Madrid"
"Y_GE15","ES30",2009,13.9,"Comunidad de Madrid"
"Y_GE15","ES4",2009,17,"Centro (ES)"
"Y_GE15","ES41",2009,14,"Castilla y León"
"Y_GE15","ES42",2009,18.9,"Castilla-la Mancha"
"Y_GE15","ES43",2009,20.6,"Extremadura"
"Y_GE15","ES5",2009,18,"Este (ES)"
"Y_GE15","ES51",2009,16.2,"Cataluña"
"Y_GE15","ES52",2009,20.8,"Comunidad Valenciana"
"Y_GE15","ES53",2009,17.9,"Illes Balears"
"Y_GE15","ES6",2009,24.4,"Sur (ES)"
"Y_GE15","ES61",2009,25.2,"Andalucía"
"Y_GE15","ES62",2009,20.3,"Región de Murcia"
"Y_GE15","ES63",2009,18.5,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2009,23.5,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2009,26,"Canarias (ES)"
"Y_GE15","ES70",2009,26,"Canarias (ES)"
"Y_GE15","EU15",2009,9,"European Union (15 countries)"
"Y_GE15","EU27",2009,8.9,"European Union (27 countries)"
"Y_GE15","EU28",2009,8.9,"European Union (28 countries)"
"Y_GE15","FI",2009,8.2,"Finland"
"Y_GE15","FI1",2009,8.3,"Manner-Suomi"
"Y_GE15","FI19",2009,9,"Länsi-Suomi"
"Y_GE15","FI1B",2009,6.2,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2009,8.1,"Etelä-Suomi"
"Y_GE15","FI1D",2009,10.5,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2009,NA,"Åland"
"Y_GE15","FI20",2009,NA,"Åland"
"Y_GE15","FR",2009,9.1,"France"
"Y_GE15","FR1",2009,8.1,"Île de France"
"Y_GE15","FR10",2009,8.1,"Île de France"
"Y_GE15","FR2",2009,8.4,"Bassin Parisien"
"Y_GE15","FR21",2009,9.2,"Champagne-Ardenne"
"Y_GE15","FR22",2009,10.3,"Picardie"
"Y_GE15","FR23",2009,10,"Haute-Normandie"
"Y_GE15","FR24",2009,6.7,"Centre (FR)"
"Y_GE15","FR25",2009,6.9,"Basse-Normandie"
"Y_GE15","FR26",2009,7.9,"Bourgogne"
"Y_GE15","FR3",2009,13.1,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2009,13.1,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2009,9.6,"Est (FR)"
"Y_GE15","FR41",2009,11.2,"Lorraine"
"Y_GE15","FR42",2009,8.2,"Alsace"
"Y_GE15","FR43",2009,8.9,"Franche-Comté"
"Y_GE15","FR5",2009,7,"Ouest (FR)"
"Y_GE15","FR51",2009,7.6,"Pays de la Loire"
"Y_GE15","FR52",2009,5.6,"Bretagne"
"Y_GE15","FR53",2009,8.4,"Poitou-Charentes"
"Y_GE15","FR6",2009,8.3,"Sud-Ouest (FR)"
"Y_GE15","FR61",2009,8.3,"Aquitaine"
"Y_GE15","FR62",2009,8.7,"Midi-Pyrénées"
"Y_GE15","FR63",2009,6.2,"Limousin"
"Y_GE15","FR7",2009,8.2,"Centre-Est (FR)"
"Y_GE15","FR71",2009,8.4,"Rhône-Alpes"
"Y_GE15","FR72",2009,7.4,"Auvergne"
"Y_GE15","FR8",2009,10.4,"Méditerranée"
"Y_GE15","FR81",2009,13.3,"Languedoc-Roussillon"
"Y_GE15","FR82",2009,9.2,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2009,NA,"Corse"
"Y_GE15","FR9",2009,24.4,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2009,23.4,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2009,21.8,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2009,20.2,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2009,27.1,"Réunion (NUTS 2010)"
"Y_GE15","HR",2009,9.2,"Croatia"
"Y_GE15","HR0",2009,9.2,"Hrvatska"
"Y_GE15","HR03",2009,9.6,"Jadranska Hrvatska"
"Y_GE15","HR04",2009,9,"Kontinentalna Hrvatska"
"Y_GE15","HU",2009,10,"Hungary"
"Y_GE15","HU1",2009,6.5,"Közép-Magyarország"
"Y_GE15","HU10",2009,6.5,"Közép-Magyarország"
"Y_GE15","HU2",2009,9.6,"Dunántúl"
"Y_GE15","HU21",2009,9.2,"Közép-Dunántúl"
"Y_GE15","HU22",2009,8.7,"Nyugat-Dunántúl"
"Y_GE15","HU23",2009,11.2,"Dél-Dunántúl"
"Y_GE15","HU3",2009,13.3,"Alföld és Észak"
"Y_GE15","HU31",2009,15.3,"Észak-Magyarország"
"Y_GE15","HU32",2009,14.1,"Észak-Alföld"
"Y_GE15","HU33",2009,10.6,"Dél-Alföld"
"Y_GE15","IE",2009,12,"Ireland"
"Y_GE15","IE0",2009,12,"Éire/Ireland"
"Y_GE15","IE01",2009,13.4,"Border, Midland and Western"
"Y_GE15","IE02",2009,11.5,"Southern and Eastern"
"Y_GE15","IS",2009,7.2,"Iceland"
"Y_GE15","IS0",2009,7.2,"Ísland"
"Y_GE15","IS00",2009,7.2,"Ísland"
"Y_GE15","IT",2009,7.7,"Italy"
"Y_GE15","ITC",2009,5.7,"Nord-Ovest"
"Y_GE15","ITC1",2009,6.8,"Piemonte"
"Y_GE15","ITC2",2009,4.5,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2009,5.8,"Liguria"
"Y_GE15","ITC4",2009,5.3,"Lombardia"
"Y_GE15","ITF",2009,11.9,"Sud"
"Y_GE15","ITF1",2009,8,"Abruzzo"
"Y_GE15","ITF2",2009,9,"Molise"
"Y_GE15","ITF3",2009,12.9,"Campania"
"Y_GE15","ITF4",2009,12.6,"Puglia"
"Y_GE15","ITF5",2009,11.2,"Basilicata"
"Y_GE15","ITF6",2009,11.3,"Calabria"
"Y_GE15","ITG",2009,13.6,"Isole"
"Y_GE15","ITG1",2009,13.8,"Sicilia"
"Y_GE15","ITG2",2009,13.2,"Sardegna"
"Y_GE15","ITH",2009,4.6,"Nord-Est"
"Y_GE15","ITH1",2009,2.9,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2009,3.5,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2009,4.7,"Veneto"
"Y_GE15","ITH4",2009,5.2,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2009,4.7,"Emilia-Romagna"
"Y_GE15","ITI",2009,7.2,"Centro (IT)"
"Y_GE15","ITI1",2009,5.8,"Toscana"
"Y_GE15","ITI2",2009,6.6,"Umbria"
"Y_GE15","ITI3",2009,6.6,"Marche"
"Y_GE15","ITI4",2009,8.4,"Lazio"
"Y_GE15","LT",2009,13.8,"Lithuania"
"Y_GE15","LT0",2009,13.8,"Lietuva"
"Y_GE15","LT00",2009,13.8,"Lietuva"
"Y_GE15","LU",2009,5.1,"Luxembourg"
"Y_GE15","LU0",2009,5.1,"Luxembourg"
"Y_GE15","LU00",2009,5.1,"Luxembourg"
"Y_GE15","LV",2009,17.5,"Latvia"
"Y_GE15","LV0",2009,17.5,"Latvija"
"Y_GE15","LV00",2009,17.5,"Latvija"
"Y_GE15","MK",2009,32.2,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2009,32.2,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2009,32.2,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2009,6.9,"Malta"
"Y_GE15","MT0",2009,6.9,"Malta"
"Y_GE15","MT00",2009,6.9,"Malta"
"Y_GE15","NL",2009,3.4,"Netherlands"
"Y_GE15","NL1",2009,4.2,"Noord-Nederland"
"Y_GE15","NL11",2009,4.8,"Groningen"
"Y_GE15","NL12",2009,3.5,"Friesland (NL)"
"Y_GE15","NL13",2009,4.2,"Drenthe"
"Y_GE15","NL2",2009,3.1,"Oost-Nederland"
"Y_GE15","NL21",2009,3.6,"Overijssel"
"Y_GE15","NL22",2009,2.8,"Gelderland"
"Y_GE15","NL23",2009,3.6,"Flevoland"
"Y_GE15","NL3",2009,3.3,"West-Nederland"
"Y_GE15","NL31",2009,2.9,"Utrecht"
"Y_GE15","NL32",2009,3.2,"Noord-Holland"
"Y_GE15","NL33",2009,3.6,"Zuid-Holland"
"Y_GE15","NL34",2009,2.1,"Zeeland"
"Y_GE15","NL4",2009,3.6,"Zuid-Nederland"
"Y_GE15","NL41",2009,3.2,"Noord-Brabant"
"Y_GE15","NL42",2009,4.4,"Limburg (NL)"
"Y_GE15","NO",2009,3.1,"Norway"
"Y_GE15","NO0",2009,3.1,"Norge"
"Y_GE15","NO01",2009,3.6,"Oslo og Akershus"
"Y_GE15","NO02",2009,2.5,"Hedmark og Oppland"
"Y_GE15","NO03",2009,3.4,"Sør-Østlandet"
"Y_GE15","NO04",2009,2.2,"Agder og Rogaland"
"Y_GE15","NO05",2009,2.4,"Vestlandet"
"Y_GE15","NO06",2009,3.7,"Trøndelag"
"Y_GE15","NO07",2009,3.7,"Nord-Norge"
"Y_GE15","PL",2009,8.2,"Poland"
"Y_GE15","PL1",2009,6.5,"Region Centralny"
"Y_GE15","PL11",2009,7.6,"Lódzkie"
"Y_GE15","PL12",2009,6,"Mazowieckie"
"Y_GE15","PL2",2009,7.2,"Region Poludniowy"
"Y_GE15","PL21",2009,7.9,"Malopolskie"
"Y_GE15","PL22",2009,6.7,"Slaskie"
"Y_GE15","PL3",2009,9.6,"Region Wschodni"
"Y_GE15","PL31",2009,9.7,"Lubelskie"
"Y_GE15","PL32",2009,10.1,"Podkarpackie"
"Y_GE15","PL33",2009,10.8,"Swietokrzyskie"
"Y_GE15","PL34",2009,7.1,"Podlaskie"
"Y_GE15","PL4",2009,8.6,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2009,7.5,"Wielkopolskie"
"Y_GE15","PL42",2009,10.4,"Zachodniopomorskie"
"Y_GE15","PL43",2009,9.6,"Lubuskie"
"Y_GE15","PL5",2009,10,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2009,10.1,"Dolnoslaskie"
"Y_GE15","PL52",2009,9.9,"Opolskie"
"Y_GE15","PL6",2009,8.5,"Region Pólnocny"
"Y_GE15","PL61",2009,10.4,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2009,8.5,"Warminsko-Mazurskie"
"Y_GE15","PL63",2009,6.4,"Pomorskie"
"Y_GE15","PT",2009,9.4,"Portugal"
"Y_GE15","PT1",2009,9.5,"Continente"
"Y_GE15","PT11",2009,10.9,"Norte"
"Y_GE15","PT15",2009,10.4,"Algarve"
"Y_GE15","PT16",2009,6.8,"Centro (PT)"
"Y_GE15","PT17",2009,9.8,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2009,10.5,"Alentejo"
"Y_GE15","PT2",2009,6.7,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2009,6.7,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2009,7.5,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2009,7.5,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2009,6.9,"Romania"
"Y_GE15","RO1",2009,8.1,"Macroregiunea unu"
"Y_GE15","RO11",2009,5.6,"Nord-Vest"
"Y_GE15","RO12",2009,10.7,"Centru"
"Y_GE15","RO2",2009,6.6,"Macroregiunea doi"
"Y_GE15","RO21",2009,6,"Nord-Est"
"Y_GE15","RO22",2009,7.5,"Sud-Est"
"Y_GE15","RO3",2009,6.4,"Macroregiunea trei"
"Y_GE15","RO31",2009,8,"Sud - Muntenia"
"Y_GE15","RO32",2009,4,"Bucuresti - Ilfov"
"Y_GE15","RO4",2009,6.5,"Macroregiunea patru"
"Y_GE15","RO41",2009,6.8,"Sud-Vest Oltenia"
"Y_GE15","RO42",2009,6,"Vest"
"Y_GE15","SE",2009,8.4,"Sweden"
"Y_GE15","SE1",2009,7.8,"Östra Sverige"
"Y_GE15","SE11",2009,6.8,"Stockholm"
"Y_GE15","SE12",2009,9.3,"Östra Mellansverige"
"Y_GE15","SE2",2009,8.5,"Södra Sverige"
"Y_GE15","SE21",2009,8.1,"Småland med öarna"
"Y_GE15","SE22",2009,8.7,"Sydsverige"
"Y_GE15","SE23",2009,8.6,"Västsverige"
"Y_GE15","SE3",2009,9.1,"Norra Sverige"
"Y_GE15","SE31",2009,9.4,"Norra Mellansverige"
"Y_GE15","SE32",2009,8.9,"Mellersta Norrland"
"Y_GE15","SE33",2009,8.9,"Övre Norrland"
"Y_GE15","SI",2009,5.9,"Slovenia"
"Y_GE15","SI0",2009,5.9,"Slovenija"
"Y_GE15","SI01",2009,6.8,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2009,4.8,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2009,12,"Slovakia"
"Y_GE15","SK0",2009,12,"Slovensko"
"Y_GE15","SK01",2009,4.6,"Bratislavský kraj"
"Y_GE15","SK02",2009,9.9,"Západné Slovensko"
"Y_GE15","SK03",2009,14.6,"Stredné Slovensko"
"Y_GE15","SK04",2009,15.9,"Východné Slovensko"
"Y_GE15","TR",2009,12.6,"Turkey"
"Y_GE15","TR1",2009,15.9,"Istanbul"
"Y_GE15","TR10",2009,15.9,"Istanbul"
"Y_GE15","TR2",2009,9.4,"Bati Marmara"
"Y_GE15","TR21",2009,11.6,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2009,7.1,"Balikesir, Çanakkale"
"Y_GE15","TR3",2009,12.9,"Ege"
"Y_GE15","TR31",2009,15.4,"Izmir"
"Y_GE15","TR32",2009,12.8,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2009,9.6,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2009,12.7,"Dogu Marmara"
"Y_GE15","TR41",2009,12.6,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2009,12.8,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2009,11.1,"Bati Anadolu"
"Y_GE15","TR51",2009,12.2,"Ankara"
"Y_GE15","TR52",2009,8.8,"Konya, Karaman"
"Y_GE15","TR6",2009,15.4,"Akdeniz"
"Y_GE15","TR61",2009,10.1,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2009,19.9,"Adana, Mersin"
"Y_GE15","TR63",2009,14.8,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2009,12.5,"Orta Anadolu"
"Y_GE15","TR71",2009,14.2,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2009,11.2,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2009,6.5,"Bati Karadeniz"
"Y_GE15","TR81",2009,6.7,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2009,8.4,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2009,6,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2009,4.2,"Dogu Karadeniz"
"Y_GE15","TR90",2009,4.2,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2009,6.9,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2009,6.3,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2009,7.5,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2009,14.7,"Ortadogu Anadolu"
"Y_GE15","TRB1",2009,14.8,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2009,14.6,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2009,15.1,"Güneydogu Anadolu"
"Y_GE15","TRC1",2009,14.3,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2009,16.7,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2009,13.8,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2009,7.5,"United Kingdom"
"Y_GE15","UKC",2009,9.1,"North East (UK)"
"Y_GE15","UKC1",2009,8.3,"Tees Valley and Durham"
"Y_GE15","UKC2",2009,9.8,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2009,8.3,"North West (UK)"
"Y_GE15","UKD1",2009,6.4,"Cumbria"
"Y_GE15","UKD3",2009,9.5,"Greater Manchester"
"Y_GE15","UKD4",2009,7.2,"Lancashire"
"Y_GE15","UKD6",2009,6,"Cheshire"
"Y_GE15","UKD7",2009,9.6,"Merseyside"
"Y_GE15","UKE",2009,8.5,"Yorkshire and The Humber"
"Y_GE15","UKE1",2009,9.4,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2009,5.4,"North Yorkshire"
"Y_GE15","UKE3",2009,9.6,"South Yorkshire"
"Y_GE15","UKE4",2009,8.6,"West Yorkshire"
"Y_GE15","UKF",2009,7.1,"East Midlands (UK)"
"Y_GE15","UKF1",2009,7.2,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2009,7.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2009,6.3,"Lincolnshire"
"Y_GE15","UKG",2009,9.6,"West Midlands (UK)"
"Y_GE15","UKG1",2009,6.4,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2009,7.1,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2009,13,"West Midlands"
"Y_GE15","UKH",2009,6.2,"East of England"
"Y_GE15","UKH1",2009,5.9,"East Anglia"
"Y_GE15","UKH2",2009,5.9,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2009,6.9,"Essex"
"Y_GE15","UKI",2009,9,"London"
"Y_GE15","UKI1",2009,9.5,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2009,8.6,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2009,5.8,"South East (UK)"
"Y_GE15","UKJ1",2009,5.4,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2009,5.6,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2009,5.2,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2009,7.3,"Kent"
"Y_GE15","UKK",2009,6.1,"South West (UK)"
"Y_GE15","UKK1",2009,5.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2009,6.5,"Dorset and Somerset"
"Y_GE15","UKK3",2009,5.1,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2009,7.1,"Devon"
"Y_GE15","UKL",2009,8,"Wales"
"Y_GE15","UKL1",2009,8.9,"West Wales and The Valleys"
"Y_GE15","UKL2",2009,6.7,"East Wales"
"Y_GE15","UKM",2009,6.9,"Scotland"
"Y_GE15","UKM2",2009,7.6,"Eastern Scotland"
"Y_GE15","UKM3",2009,7.5,"South Western Scotland"
"Y_GE15","UKM5",2009,3.6,"North Eastern Scotland"
"Y_GE15","UKM6",2009,4.3,"Highlands and Islands"
"Y_GE15","UKN",2009,6.4,"Northern Ireland (UK)"
"Y_GE15","UKN0",2009,6.4,"Northern Ireland (UK)"
"Y_GE25","AT",2009,4.4,"Austria"
"Y_GE25","AT1",2009,5.6,"Ostösterreich"
"Y_GE25","AT11",2009,4.4,"Burgenland (AT)"
"Y_GE25","AT12",2009,3.6,"Niederösterreich"
"Y_GE25","AT13",2009,7.7,"Wien"
"Y_GE25","AT2",2009,4,"Südösterreich"
"Y_GE25","AT21",2009,3.8,"Kärnten"
"Y_GE25","AT22",2009,4,"Steiermark"
"Y_GE25","AT3",2009,3.3,"Westösterreich"
"Y_GE25","AT31",2009,3.6,"Oberösterreich"
"Y_GE25","AT32",2009,2.8,"Salzburg"
"Y_GE25","AT33",2009,2.6,"Tirol"
"Y_GE25","AT34",2009,4.5,"Vorarlberg"
"Y_GE25","BE",2009,6.5,"Belgium"
"Y_GE25","BE1",2009,14.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2009,14.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2009,3.9,"Vlaams Gewest"
"Y_GE25","BE21",2009,4.8,"Prov. Antwerpen"
"Y_GE25","BE22",2009,4,"Prov. Limburg (BE)"
"Y_GE25","BE23",2009,3.3,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2009,3.8,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2009,3.4,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2009,9.1,"Région wallonne"
"Y_GE25","BE31",2009,6,"Prov. Brabant Wallon"
"Y_GE25","BE32",2009,10.4,"Prov. Hainaut"
"Y_GE25","BE33",2009,10.2,"Prov. Liège"
"Y_GE25","BE34",2009,5.7,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2009,8.1,"Prov. Namur"
"Y_GE25","BG",2009,6,"Bulgaria"
"Y_GE25","BG3",2009,7.3,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2009,7.5,"Severozapaden"
"Y_GE25","BG32",2009,7.1,"Severen tsentralen"
"Y_GE25","BG33",2009,9.3,"Severoiztochen"
"Y_GE25","BG34",2009,5.6,"Yugoiztochen"
"Y_GE25","BG4",2009,4.7,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2009,3.6,"Yugozapaden"
"Y_GE25","BG42",2009,6.4,"Yuzhen tsentralen"
"Y_GE25","CH",2009,3.4,"Switzerland"
"Y_GE25","CH0",2009,3.4,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2009,4.7,"Région lémanique"
"Y_GE25","CH02",2009,2.9,"Espace Mittelland"
"Y_GE25","CH03",2009,3.8,"Nordwestschweiz"
"Y_GE25","CH04",2009,3.2,"Zürich"
"Y_GE25","CH05",2009,3.2,"Ostschweiz"
"Y_GE25","CH06",2009,2.2,"Zentralschweiz"
"Y_GE25","CH07",2009,4,"Ticino"
"Y_GE25","CY",2009,4.4,"Cyprus"
"Y_GE25","CY0",2009,4.4,"Kypros"
"Y_GE25","CY00",2009,4.4,"Kypros"
"Y_GE25","CZ",2009,5.8,"Czech Republic"
"Y_GE25","CZ0",2009,5.8,"Ceská republika"
"Y_GE25","CZ01",2009,2.6,"Praha"
"Y_GE25","CZ02",2009,3.4,"Strední Cechy"
"Y_GE25","CZ03",2009,4.5,"Jihozápad"
"Y_GE25","CZ04",2009,8.9,"Severozápad"
"Y_GE25","CZ05",2009,6.6,"Severovýchod"
"Y_GE25","CZ06",2009,5.7,"Jihovýchod"
"Y_GE25","CZ07",2009,6.6,"Strední Morava"
"Y_GE25","CZ08",2009,8.6,"Moravskoslezsko"
"Y_GE25","DE",2009,7.3,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2009,4.7,"Baden-Württemberg"
"Y_GE25","DE11",2009,4.7,"Stuttgart"
"Y_GE25","DE12",2009,5.1,"Karlsruhe"
"Y_GE25","DE13",2009,4.1,"Freiburg"
"Y_GE25","DE14",2009,4.9,"Tübingen"
"Y_GE25","DE2",2009,4.7,"Bayern"
"Y_GE25","DE21",2009,4,"Oberbayern"
"Y_GE25","DE22",2009,4.7,"Niederbayern"
"Y_GE25","DE23",2009,4.6,"Oberpfalz"
"Y_GE25","DE24",2009,5.7,"Oberfranken"
"Y_GE25","DE25",2009,6,"Mittelfranken"
"Y_GE25","DE26",2009,5.1,"Unterfranken"
"Y_GE25","DE27",2009,4.3,"Schwaben"
"Y_GE25","DE3",2009,13.3,"Berlin"
"Y_GE25","DE30",2009,13.3,"Berlin"
"Y_GE25","DE4",2009,10.6,"Brandenburg"
"Y_GE25","DE40",2009,10.6,"Brandenburg"
"Y_GE25","DE5",2009,9.4,"Bremen"
"Y_GE25","DE50",2009,9.4,"Bremen"
"Y_GE25","DE6",2009,6.8,"Hamburg"
"Y_GE25","DE60",2009,6.8,"Hamburg"
"Y_GE25","DE7",2009,5.8,"Hessen"
"Y_GE25","DE71",2009,5.8,"Darmstadt"
"Y_GE25","DE72",2009,5.8,"Gießen"
"Y_GE25","DE73",2009,6,"Kassel"
"Y_GE25","DE8",2009,13.7,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2009,13.7,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2009,6.5,"Niedersachsen"
"Y_GE25","DE91",2009,8.2,"Braunschweig"
"Y_GE25","DE92",2009,7.5,"Hannover"
"Y_GE25","DE93",2009,4.9,"Lüneburg"
"Y_GE25","DE94",2009,5.4,"Weser-Ems"
"Y_GE25","DEA",2009,7.3,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2009,7.1,"Düsseldorf"
"Y_GE25","DEA2",2009,6.7,"Köln"
"Y_GE25","DEA3",2009,6.9,"Münster"
"Y_GE25","DEA4",2009,7.2,"Detmold"
"Y_GE25","DEA5",2009,8.6,"Arnsberg"
"Y_GE25","DEB",2009,5.3,"Rheinland-Pfalz"
"Y_GE25","DEB1",2009,6.1,"Koblenz"
"Y_GE25","DEB2",2009,4.1,"Trier"
"Y_GE25","DEB3",2009,5.1,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2009,7.6,"Saarland"
"Y_GE25","DEC0",2009,7.6,"Saarland"
"Y_GE25","DED",2009,12.1,"Sachsen"
"Y_GE25","DED2",2009,11.4,"Dresden"
"Y_GE25","DED4",2009,12.5,"Chemnitz"
"Y_GE25","DED5",2009,12.8,"Leipzig"
"Y_GE25","DEE",2009,13.4,"Sachsen-Anhalt"
"Y_GE25","DEE0",2009,13.4,"Sachsen-Anhalt"
"Y_GE25","DEF",2009,6.9,"Schleswig-Holstein"
"Y_GE25","DEF0",2009,6.9,"Schleswig-Holstein"
"Y_GE25","DEG",2009,10.5,"Thüringen"
"Y_GE25","DEG0",2009,10.5,"Thüringen"
"Y_GE25","DK",2009,4.9,"Denmark"
"Y_GE25","DK0",2009,4.9,"Danmark"
"Y_GE25","DK01",2009,5.1,"Hovedstaden"
"Y_GE25","DK02",2009,4.1,"Sjælland"
"Y_GE25","DK03",2009,4.8,"Syddanmark"
"Y_GE25","DK04",2009,4.8,"Midtjylland"
"Y_GE25","DK05",2009,6,"Nordjylland"
"Y_GE25","EA17",2009,8.2,"Euro area (17 countries)"
"Y_GE25","EA18",2009,8.3,"Euro area (18 countries)"
"Y_GE25","EA19",2009,8.3,"Euro area (19 countries)"
"Y_GE25","EE",2009,11.9,"Estonia"
"Y_GE25","EE0",2009,11.9,"Eesti"
"Y_GE25","EE00",2009,11.9,"Eesti"
"Y_GE25","EL",2009,8.3,"Greece"
"Y_GE25","EL1",2009,8.9,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2009,9.4,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2009,8.8,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2009,11.1,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2009,7.9,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2009,7.9,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2009,9.2,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2009,7.9,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2009,7.7,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2009,8.5,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2009,6.8,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2009,8.1,"Attiki"
"Y_GE25","EL30",2009,8.1,"Attiki"
"Y_GE25","EL4",2009,8.4,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2009,5.2,"Voreio Aigaio"
"Y_GE25","EL42",2009,11,"Notio Aigaio"
"Y_GE25","EL43",2009,7.9,"Kriti"
"Y_GE25","ES",2009,15.7,"Spain"
"Y_GE25","ES1",2009,11,"Noroeste (ES)"
"Y_GE25","ES11",2009,10.9,"Galicia"
"Y_GE25","ES12",2009,11.6,"Principado de Asturias"
"Y_GE25","ES13",2009,10.5,"Cantabria"
"Y_GE25","ES2",2009,10.2,"Noreste (ES)"
"Y_GE25","ES21",2009,9.8,"País Vasco"
"Y_GE25","ES22",2009,9,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2009,10.6,"La Rioja"
"Y_GE25","ES24",2009,11.3,"Aragón"
"Y_GE25","ES3",2009,11.9,"Comunidad de Madrid"
"Y_GE25","ES30",2009,11.9,"Comunidad de Madrid"
"Y_GE25","ES4",2009,14.9,"Centro (ES)"
"Y_GE25","ES41",2009,12.3,"Castilla y León"
"Y_GE25","ES42",2009,16.6,"Castilla-la Mancha"
"Y_GE25","ES43",2009,18,"Extremadura"
"Y_GE25","ES5",2009,15.9,"Este (ES)"
"Y_GE25","ES51",2009,14.1,"Cataluña"
"Y_GE25","ES52",2009,18.6,"Comunidad Valenciana"
"Y_GE25","ES53",2009,16.3,"Illes Balears"
"Y_GE25","ES6",2009,22.1,"Sur (ES)"
"Y_GE25","ES61",2009,22.7,"Andalucía"
"Y_GE25","ES62",2009,18.7,"Región de Murcia"
"Y_GE25","ES63",2009,16.4,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2009,21.8,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2009,23.7,"Canarias (ES)"
"Y_GE25","ES70",2009,23.7,"Canarias (ES)"
"Y_GE25","EU15",2009,7.7,"European Union (15 countries)"
"Y_GE25","EU27",2009,7.6,"European Union (27 countries)"
"Y_GE25","EU28",2009,7.6,"European Union (28 countries)"
"Y_GE25","FI",2009,6.4,"Finland"
"Y_GE25","FI1",2009,6.4,"Manner-Suomi"
"Y_GE25","FI19",2009,7.2,"Länsi-Suomi"
"Y_GE25","FI1B",2009,4.6,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2009,6.2,"Etelä-Suomi"
"Y_GE25","FI1D",2009,8.4,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2009,NA,"Åland"
"Y_GE25","FI20",2009,NA,"Åland"
"Y_GE25","FR",2009,7.4,"France"
"Y_GE25","FR1",2009,6.8,"Île de France"
"Y_GE25","FR10",2009,6.8,"Île de France"
"Y_GE25","FR2",2009,6.6,"Bassin Parisien"
"Y_GE25","FR21",2009,7.8,"Champagne-Ardenne"
"Y_GE25","FR22",2009,8.2,"Picardie"
"Y_GE25","FR23",2009,7.9,"Haute-Normandie"
"Y_GE25","FR24",2009,5.3,"Centre (FR)"
"Y_GE25","FR25",2009,5.3,"Basse-Normandie"
"Y_GE25","FR26",2009,5.9,"Bourgogne"
"Y_GE25","FR3",2009,9.9,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2009,9.9,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2009,7.9,"Est (FR)"
"Y_GE25","FR41",2009,9.1,"Lorraine"
"Y_GE25","FR42",2009,6.8,"Alsace"
"Y_GE25","FR43",2009,7.3,"Franche-Comté"
"Y_GE25","FR5",2009,5.7,"Ouest (FR)"
"Y_GE25","FR51",2009,6.2,"Pays de la Loire"
"Y_GE25","FR52",2009,4.6,"Bretagne"
"Y_GE25","FR53",2009,6.8,"Poitou-Charentes"
"Y_GE25","FR6",2009,6.8,"Sud-Ouest (FR)"
"Y_GE25","FR61",2009,6.9,"Aquitaine"
"Y_GE25","FR62",2009,7.3,"Midi-Pyrénées"
"Y_GE25","FR63",2009,5.1,"Limousin"
"Y_GE25","FR7",2009,6.6,"Centre-Est (FR)"
"Y_GE25","FR71",2009,6.6,"Rhône-Alpes"
"Y_GE25","FR72",2009,6.4,"Auvergne"
"Y_GE25","FR8",2009,8.4,"Méditerranée"
"Y_GE25","FR81",2009,10.7,"Languedoc-Roussillon"
"Y_GE25","FR82",2009,7.4,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2009,NA,"Corse"
"Y_GE25","FR9",2009,21.2,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2009,20.6,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2009,18.7,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2009,17.8,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2009,23.7,"Réunion (NUTS 2010)"
"Y_GE25","HR",2009,7.5,"Croatia"
"Y_GE25","HR0",2009,7.5,"Hrvatska"
"Y_GE25","HR03",2009,8.3,"Jadranska Hrvatska"
"Y_GE25","HR04",2009,7.1,"Kontinentalna Hrvatska"
"Y_GE25","HU",2009,8.8,"Hungary"
"Y_GE25","HU1",2009,5.8,"Közép-Magyarország"
"Y_GE25","HU10",2009,5.8,"Közép-Magyarország"
"Y_GE25","HU2",2009,8.3,"Dunántúl"
"Y_GE25","HU21",2009,8.1,"Közép-Dunántúl"
"Y_GE25","HU22",2009,7.5,"Nyugat-Dunántúl"
"Y_GE25","HU23",2009,9.4,"Dél-Dunántúl"
"Y_GE25","HU3",2009,11.7,"Alföld és Észak"
"Y_GE25","HU31",2009,13.5,"Észak-Magyarország"
"Y_GE25","HU32",2009,12.4,"Észak-Alföld"
"Y_GE25","HU33",2009,9.4,"Dél-Alföld"
"Y_GE25","IE",2009,10.1,"Ireland"
"Y_GE25","IE0",2009,10.1,"Éire/Ireland"
"Y_GE25","IE01",2009,11.1,"Border, Midland and Western"
"Y_GE25","IE02",2009,9.7,"Southern and Eastern"
"Y_GE25","IS",2009,5.5,"Iceland"
"Y_GE25","IS0",2009,5.5,"Ísland"
"Y_GE25","IS00",2009,5.5,"Ísland"
"Y_GE25","IT",2009,6.4,"Italy"
"Y_GE25","ITC",2009,4.7,"Nord-Ovest"
"Y_GE25","ITC1",2009,5.6,"Piemonte"
"Y_GE25","ITC2",2009,3.6,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2009,5.1,"Liguria"
"Y_GE25","ITC4",2009,4.3,"Lombardia"
"Y_GE25","ITF",2009,9.9,"Sud"
"Y_GE25","ITF1",2009,6.9,"Abruzzo"
"Y_GE25","ITF2",2009,7.7,"Molise"
"Y_GE25","ITF3",2009,10.6,"Campania"
"Y_GE25","ITF4",2009,10.5,"Puglia"
"Y_GE25","ITF5",2009,9.1,"Basilicata"
"Y_GE25","ITF6",2009,9.6,"Calabria"
"Y_GE25","ITG",2009,11.3,"Isole"
"Y_GE25","ITG1",2009,11.5,"Sicilia"
"Y_GE25","ITG2",2009,10.8,"Sardegna"
"Y_GE25","ITH",2009,3.9,"Nord-Est"
"Y_GE25","ITH1",2009,2.2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2009,2.9,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2009,4,"Veneto"
"Y_GE25","ITH4",2009,4.4,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2009,3.9,"Emilia-Romagna"
"Y_GE25","ITI",2009,6,"Centro (IT)"
"Y_GE25","ITI1",2009,5,"Toscana"
"Y_GE25","ITI2",2009,5.7,"Umbria"
"Y_GE25","ITI3",2009,5.4,"Marche"
"Y_GE25","ITI4",2009,6.9,"Lazio"
"Y_GE25","LT",2009,12.2,"Lithuania"
"Y_GE25","LT0",2009,12.2,"Lietuva"
"Y_GE25","LT00",2009,12.2,"Lietuva"
"Y_GE25","LU",2009,4.1,"Luxembourg"
"Y_GE25","LU0",2009,4.1,"Luxembourg"
"Y_GE25","LU00",2009,4.1,"Luxembourg"
"Y_GE25","LV",2009,15.4,"Latvia"
"Y_GE25","LV0",2009,15.4,"Latvija"
"Y_GE25","LV00",2009,15.4,"Latvija"
"Y_GE25","MK",2009,29,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2009,29,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2009,29,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2009,5.3,"Malta"
"Y_GE25","MT0",2009,5.3,"Malta"
"Y_GE25","MT00",2009,5.3,"Malta"
"Y_GE25","NL",2009,2.8,"Netherlands"
"Y_GE25","NL1",2009,3.4,"Noord-Nederland"
"Y_GE25","NL11",2009,3.9,"Groningen"
"Y_GE25","NL12",2009,2.8,"Friesland (NL)"
"Y_GE25","NL13",2009,3.7,"Drenthe"
"Y_GE25","NL2",2009,2.6,"Oost-Nederland"
"Y_GE25","NL21",2009,3.2,"Overijssel"
"Y_GE25","NL22",2009,2.2,"Gelderland"
"Y_GE25","NL23",2009,2.6,"Flevoland"
"Y_GE25","NL3",2009,2.7,"West-Nederland"
"Y_GE25","NL31",2009,2.3,"Utrecht"
"Y_GE25","NL32",2009,2.7,"Noord-Holland"
"Y_GE25","NL33",2009,2.8,"Zuid-Holland"
"Y_GE25","NL34",2009,1.8,"Zeeland"
"Y_GE25","NL4",2009,2.9,"Zuid-Nederland"
"Y_GE25","NL41",2009,2.6,"Noord-Brabant"
"Y_GE25","NL42",2009,3.6,"Limburg (NL)"
"Y_GE25","NO",2009,2.1,"Norway"
"Y_GE25","NO0",2009,2.1,"Norge"
"Y_GE25","NO01",2009,2.7,"Oslo og Akershus"
"Y_GE25","NO02",2009,1.6,"Hedmark og Oppland"
"Y_GE25","NO03",2009,2.3,"Sør-Østlandet"
"Y_GE25","NO04",2009,1.7,"Agder og Rogaland"
"Y_GE25","NO05",2009,1.5,"Vestlandet"
"Y_GE25","NO06",2009,2.6,"Trøndelag"
"Y_GE25","NO07",2009,2.1,"Nord-Norge"
"Y_GE25","PL",2009,6.8,"Poland"
"Y_GE25","PL1",2009,5.5,"Region Centralny"
"Y_GE25","PL11",2009,6.5,"Lódzkie"
"Y_GE25","PL12",2009,5,"Mazowieckie"
"Y_GE25","PL2",2009,5.7,"Region Poludniowy"
"Y_GE25","PL21",2009,6,"Malopolskie"
"Y_GE25","PL22",2009,5.5,"Slaskie"
"Y_GE25","PL3",2009,7.8,"Region Wschodni"
"Y_GE25","PL31",2009,8,"Lubelskie"
"Y_GE25","PL32",2009,7.7,"Podkarpackie"
"Y_GE25","PL33",2009,9.3,"Swietokrzyskie"
"Y_GE25","PL34",2009,5.9,"Podlaskie"
"Y_GE25","PL4",2009,7.2,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2009,6,"Wielkopolskie"
"Y_GE25","PL42",2009,8.9,"Zachodniopomorskie"
"Y_GE25","PL43",2009,8.2,"Lubuskie"
"Y_GE25","PL5",2009,8.5,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2009,8.4,"Dolnoslaskie"
"Y_GE25","PL52",2009,8.6,"Opolskie"
"Y_GE25","PL6",2009,7.2,"Region Pólnocny"
"Y_GE25","PL61",2009,9,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2009,7.4,"Warminsko-Mazurskie"
"Y_GE25","PL63",2009,5.3,"Pomorskie"
"Y_GE25","PT",2009,8.4,"Portugal"
"Y_GE25","PT1",2009,8.6,"Continente"
"Y_GE25","PT11",2009,9.8,"Norte"
"Y_GE25","PT15",2009,9.1,"Algarve"
"Y_GE25","PT16",2009,6,"Centro (PT)"
"Y_GE25","PT17",2009,9.1,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2009,9.4,"Alentejo"
"Y_GE25","PT2",2009,5.3,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2009,5.3,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2009,6.3,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2009,6.3,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2009,5.4,"Romania"
"Y_GE25","RO1",2009,6.5,"Macroregiunea unu"
"Y_GE25","RO11",2009,4.5,"Nord-Vest"
"Y_GE25","RO12",2009,8.5,"Centru"
"Y_GE25","RO2",2009,5.3,"Macroregiunea doi"
"Y_GE25","RO21",2009,4.8,"Nord-Est"
"Y_GE25","RO22",2009,5.9,"Sud-Est"
"Y_GE25","RO3",2009,4.8,"Macroregiunea trei"
"Y_GE25","RO31",2009,6.1,"Sud - Muntenia"
"Y_GE25","RO32",2009,3,"Bucuresti - Ilfov"
"Y_GE25","RO4",2009,5.2,"Macroregiunea patru"
"Y_GE25","RO41",2009,5.5,"Sud-Vest Oltenia"
"Y_GE25","RO42",2009,4.8,"Vest"
"Y_GE25","SE",2009,5.9,"Sweden"
"Y_GE25","SE1",2009,5.6,"Östra Sverige"
"Y_GE25","SE11",2009,4.9,"Stockholm"
"Y_GE25","SE12",2009,6.6,"Östra Mellansverige"
"Y_GE25","SE2",2009,6,"Södra Sverige"
"Y_GE25","SE21",2009,5.3,"Småland med öarna"
"Y_GE25","SE22",2009,6.1,"Sydsverige"
"Y_GE25","SE23",2009,6.1,"Västsverige"
"Y_GE25","SE3",2009,6.5,"Norra Sverige"
"Y_GE25","SE31",2009,6.8,"Norra Mellansverige"
"Y_GE25","SE32",2009,5.8,"Mellersta Norrland"
"Y_GE25","SE33",2009,6.4,"Övre Norrland"
"Y_GE25","SI",2009,5,"Slovenia"
"Y_GE25","SI0",2009,5,"Slovenija"
"Y_GE25","SI01",2009,5.9,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2009,4.1,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2009,10.4,"Slovakia"
"Y_GE25","SK0",2009,10.4,"Slovensko"
"Y_GE25","SK01",2009,4.2,"Bratislavský kraj"
"Y_GE25","SK02",2009,8.6,"Západné Slovensko"
"Y_GE25","SK03",2009,12.7,"Stredné Slovensko"
"Y_GE25","SK04",2009,13.7,"Východné Slovensko"
"Y_GE25","TR",2009,10.4,"Turkey"
"Y_GE25","TR1",2009,13.7,"Istanbul"
"Y_GE25","TR10",2009,13.7,"Istanbul"
"Y_GE25","TR2",2009,7.4,"Bati Marmara"
"Y_GE25","TR21",2009,8.9,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2009,5.8,"Balikesir, Çanakkale"
"Y_GE25","TR3",2009,10.6,"Ege"
"Y_GE25","TR31",2009,12.4,"Izmir"
"Y_GE25","TR32",2009,10.9,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2009,7.5,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2009,10.5,"Dogu Marmara"
"Y_GE25","TR41",2009,10.7,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2009,10.4,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2009,9,"Bati Anadolu"
"Y_GE25","TR51",2009,9.9,"Ankara"
"Y_GE25","TR52",2009,7.2,"Konya, Karaman"
"Y_GE25","TR6",2009,13,"Akdeniz"
"Y_GE25","TR61",2009,8.4,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2009,16.8,"Adana, Mersin"
"Y_GE25","TR63",2009,13,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2009,9.9,"Orta Anadolu"
"Y_GE25","TR71",2009,11.3,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2009,9,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2009,5.2,"Bati Karadeniz"
"Y_GE25","TR81",2009,4.7,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2009,6.6,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2009,5.1,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2009,3,"Dogu Karadeniz"
"Y_GE25","TR90",2009,3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2009,5.3,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2009,4.9,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2009,5.8,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2009,11.9,"Ortadogu Anadolu"
"Y_GE25","TRB1",2009,11.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2009,12.2,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2009,12.9,"Güneydogu Anadolu"
"Y_GE25","TRC1",2009,12.2,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2009,14.7,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2009,11.2,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2009,5.6,"United Kingdom"
"Y_GE25","UKC",2009,6.5,"North East (UK)"
"Y_GE25","UKC1",2009,5.8,"Tees Valley and Durham"
"Y_GE25","UKC2",2009,7,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2009,6,"North West (UK)"
"Y_GE25","UKD1",2009,3.9,"Cumbria"
"Y_GE25","UKD3",2009,7.1,"Greater Manchester"
"Y_GE25","UKD4",2009,5.4,"Lancashire"
"Y_GE25","UKD6",2009,3.9,"Cheshire"
"Y_GE25","UKD7",2009,6.8,"Merseyside"
"Y_GE25","UKE",2009,6.2,"Yorkshire and The Humber"
"Y_GE25","UKE1",2009,6.6,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2009,4.1,"North Yorkshire"
"Y_GE25","UKE3",2009,7,"South Yorkshire"
"Y_GE25","UKE4",2009,6.5,"West Yorkshire"
"Y_GE25","UKF",2009,5.3,"East Midlands (UK)"
"Y_GE25","UKF1",2009,5.8,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2009,5.5,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2009,3.4,"Lincolnshire"
"Y_GE25","UKG",2009,7.2,"West Midlands (UK)"
"Y_GE25","UKG1",2009,4.4,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2009,5.3,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2009,9.9,"West Midlands"
"Y_GE25","UKH",2009,4.4,"East of England"
"Y_GE25","UKH1",2009,3.9,"East Anglia"
"Y_GE25","UKH2",2009,4.2,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2009,5.3,"Essex"
"Y_GE25","UKI",2009,6.9,"London"
"Y_GE25","UKI1",2009,7.4,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2009,6.6,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2009,4.1,"South East (UK)"
"Y_GE25","UKJ1",2009,3.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2009,4.2,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2009,3.7,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2009,4.7,"Kent"
"Y_GE25","UKK",2009,4.6,"South West (UK)"
"Y_GE25","UKK1",2009,4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2009,5.5,"Dorset and Somerset"
"Y_GE25","UKK3",2009,4,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2009,4.9,"Devon"
"Y_GE25","UKL",2009,5.9,"Wales"
"Y_GE25","UKL1",2009,6.3,"West Wales and The Valleys"
"Y_GE25","UKL2",2009,5.2,"East Wales"
"Y_GE25","UKM",2009,5.1,"Scotland"
"Y_GE25","UKM2",2009,5.3,"Eastern Scotland"
"Y_GE25","UKM3",2009,5.9,"South Western Scotland"
"Y_GE25","UKM5",2009,2.6,"North Eastern Scotland"
"Y_GE25","UKM6",2009,3.4,"Highlands and Islands"
"Y_GE25","UKN",2009,4.7,"Northern Ireland (UK)"
"Y_GE25","UKN0",2009,4.7,"Northern Ireland (UK)"
"Y15-24","AT",2008,8.5,"Austria"
"Y15-24","AT1",2008,11.7,"Ostösterreich"
"Y15-24","AT11",2008,NA,"Burgenland (AT)"
"Y15-24","AT12",2008,8.9,"Niederösterreich"
"Y15-24","AT13",2008,15.2,"Wien"
"Y15-24","AT2",2008,7.2,"Südösterreich"
"Y15-24","AT21",2008,NA,"Kärnten"
"Y15-24","AT22",2008,7.2,"Steiermark"
"Y15-24","AT3",2008,6.2,"Westösterreich"
"Y15-24","AT31",2008,5.4,"Oberösterreich"
"Y15-24","AT32",2008,NA,"Salzburg"
"Y15-24","AT33",2008,6.2,"Tirol"
"Y15-24","AT34",2008,NA,"Vorarlberg"
"Y15-24","BE",2008,18,"Belgium"
"Y15-24","BE1",2008,33.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2008,33.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2008,10.5,"Vlaams Gewest"
"Y15-24","BE21",2008,10.2,"Prov. Antwerpen"
"Y15-24","BE22",2008,11.7,"Prov. Limburg (BE)"
"Y15-24","BE23",2008,11.4,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2008,12,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2008,8,"Prov. West-Vlaanderen"
"Y15-24","BE3",2008,27.5,"Région wallonne"
"Y15-24","BE31",2008,19.7,"Prov. Brabant Wallon"
"Y15-24","BE32",2008,32.8,"Prov. Hainaut"
"Y15-24","BE33",2008,26.9,"Prov. Liège"
"Y15-24","BE34",2008,22.9,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2008,23.8,"Prov. Namur"
"Y15-24","BG",2008,12.7,"Bulgaria"
"Y15-24","BG3",2008,17.4,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2008,18.3,"Severozapaden"
"Y15-24","BG32",2008,17.9,"Severen tsentralen"
"Y15-24","BG33",2008,19,"Severoiztochen"
"Y15-24","BG34",2008,14.8,"Yugoiztochen"
"Y15-24","BG4",2008,7.8,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2008,6.7,"Yugozapaden"
"Y15-24","BG42",2008,9.7,"Yuzhen tsentralen"
"Y15-24","CH",2008,7,"Switzerland"
"Y15-24","CH0",2008,7,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2008,11.1,"Région lémanique"
"Y15-24","CH02",2008,7,"Espace Mittelland"
"Y15-24","CH03",2008,7.4,"Nordwestschweiz"
"Y15-24","CH04",2008,6.2,"Zürich"
"Y15-24","CH05",2008,5.1,"Ostschweiz"
"Y15-24","CH06",2008,NA,"Zentralschweiz"
"Y15-24","CH07",2008,11.2,"Ticino"
"Y15-24","CY",2008,9,"Cyprus"
"Y15-24","CY0",2008,9,"Kypros"
"Y15-24","CY00",2008,9,"Kypros"
"Y15-24","CZ",2008,9.9,"Czech Republic"
"Y15-24","CZ0",2008,9.9,"Ceská republika"
"Y15-24","CZ01",2008,4.8,"Praha"
"Y15-24","CZ02",2008,6.1,"Strední Cechy"
"Y15-24","CZ03",2008,6.6,"Jihozápad"
"Y15-24","CZ04",2008,18.2,"Severozápad"
"Y15-24","CZ05",2008,8.3,"Severovýchod"
"Y15-24","CZ06",2008,7.8,"Jihovýchod"
"Y15-24","CZ07",2008,11.2,"Strední Morava"
"Y15-24","CZ08",2008,15,"Moravskoslezsko"
"Y15-24","DE",2008,10.6,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2008,6.6,"Baden-Württemberg"
"Y15-24","DE11",2008,6.9,"Stuttgart"
"Y15-24","DE12",2008,6.5,"Karlsruhe"
"Y15-24","DE13",2008,6.3,"Freiburg"
"Y15-24","DE14",2008,6.7,"Tübingen"
"Y15-24","DE2",2008,6.1,"Bayern"
"Y15-24","DE21",2008,5,"Oberbayern"
"Y15-24","DE22",2008,NA,"Niederbayern"
"Y15-24","DE23",2008,NA,"Oberpfalz"
"Y15-24","DE24",2008,8.6,"Oberfranken"
"Y15-24","DE25",2008,7.3,"Mittelfranken"
"Y15-24","DE26",2008,6.8,"Unterfranken"
"Y15-24","DE27",2008,6.3,"Schwaben"
"Y15-24","DE3",2008,17.9,"Berlin"
"Y15-24","DE30",2008,17.9,"Berlin"
"Y15-24","DE4",2008,14.6,"Brandenburg"
"Y15-24","DE40",2008,14.6,"Brandenburg"
"Y15-24","DE5",2008,NA,"Bremen"
"Y15-24","DE50",2008,NA,"Bremen"
"Y15-24","DE6",2008,12.2,"Hamburg"
"Y15-24","DE60",2008,12.2,"Hamburg"
"Y15-24","DE7",2008,10.6,"Hessen"
"Y15-24","DE71",2008,10.1,"Darmstadt"
"Y15-24","DE72",2008,12.4,"Gießen"
"Y15-24","DE73",2008,10.3,"Kassel"
"Y15-24","DE8",2008,15,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2008,15,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2008,10.5,"Niedersachsen"
"Y15-24","DE91",2008,11.3,"Braunschweig"
"Y15-24","DE92",2008,11,"Hannover"
"Y15-24","DE93",2008,11.3,"Lüneburg"
"Y15-24","DE94",2008,9.2,"Weser-Ems"
"Y15-24","DEA",2008,11.5,"Nordrhein-Westfalen"
"Y15-24","DEA1",2008,12.7,"Düsseldorf"
"Y15-24","DEA2",2008,10.8,"Köln"
"Y15-24","DEA3",2008,8.8,"Münster"
"Y15-24","DEA4",2008,11.9,"Detmold"
"Y15-24","DEA5",2008,12.1,"Arnsberg"
"Y15-24","DEB",2008,9.7,"Rheinland-Pfalz"
"Y15-24","DEB1",2008,9.7,"Koblenz"
"Y15-24","DEB2",2008,NA,"Trier"
"Y15-24","DEB3",2008,9.8,"Rheinhessen-Pfalz"
"Y15-24","DEC",2008,14,"Saarland"
"Y15-24","DEC0",2008,14,"Saarland"
"Y15-24","DED",2008,15.7,"Sachsen"
"Y15-24","DED2",2008,17.8,"Dresden"
"Y15-24","DED4",2008,12.3,"Chemnitz"
"Y15-24","DED5",2008,16.8,"Leipzig"
"Y15-24","DEE",2008,18.2,"Sachsen-Anhalt"
"Y15-24","DEE0",2008,18.2,"Sachsen-Anhalt"
"Y15-24","DEF",2008,11.3,"Schleswig-Holstein"
"Y15-24","DEF0",2008,11.3,"Schleswig-Holstein"
"Y15-24","DEG",2008,11.8,"Thüringen"
"Y15-24","DEG0",2008,11.8,"Thüringen"
"Y15-24","DK",2008,8,"Denmark"
"Y15-24","DK0",2008,8,"Danmark"
"Y15-24","DK01",2008,7.2,"Hovedstaden"
"Y15-24","DK02",2008,9.4,"Sjælland"
"Y15-24","DK03",2008,8,"Syddanmark"
"Y15-24","DK04",2008,8.7,"Midtjylland"
"Y15-24","DK05",2008,7.4,"Nordjylland"
"Y15-24","EA17",2008,15.7,"Euro area (17 countries)"
"Y15-24","EA18",2008,15.7,"Euro area (18 countries)"
"Y15-24","EA19",2008,15.7,"Euro area (19 countries)"
"Y15-24","EE",2008,12,"Estonia"
"Y15-24","EE0",2008,12,"Eesti"
"Y15-24","EE00",2008,12,"Eesti"
"Y15-24","EL",2008,21.9,"Greece"
"Y15-24","EL1",2008,23.4,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2008,21.4,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2008,22.4,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2008,36.6,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2008,23.7,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2008,28.5,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2008,31.2,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2008,27.1,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2008,31.3,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2008,27.7,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2008,23.1,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2008,19.1,"Attiki"
"Y15-24","EL30",2008,19.1,"Attiki"
"Y15-24","EL4",2008,15,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2008,NA,"Voreio Aigaio"
"Y15-24","EL42",2008,14.9,"Notio Aigaio"
"Y15-24","EL43",2008,14,"Kriti"
"Y15-24","ES",2008,24.5,"Spain"
"Y15-24","ES1",2008,20.9,"Noroeste (ES)"
"Y15-24","ES11",2008,21.1,"Galicia"
"Y15-24","ES12",2008,21.6,"Principado de Asturias"
"Y15-24","ES13",2008,19.2,"Cantabria"
"Y15-24","ES2",2008,19.7,"Noreste (ES)"
"Y15-24","ES21",2008,19.5,"País Vasco"
"Y15-24","ES22",2008,18.8,"Comunidad Foral de Navarra"
"Y15-24","ES23",2008,21.7,"La Rioja"
"Y15-24","ES24",2008,19.8,"Aragón"
"Y15-24","ES3",2008,20.8,"Comunidad de Madrid"
"Y15-24","ES30",2008,20.8,"Comunidad de Madrid"
"Y15-24","ES4",2008,24,"Centro (ES)"
"Y15-24","ES41",2008,22.5,"Castilla y León"
"Y15-24","ES42",2008,22.9,"Castilla-la Mancha"
"Y15-24","ES43",2008,29,"Extremadura"
"Y15-24","ES5",2008,22.8,"Este (ES)"
"Y15-24","ES51",2008,20.1,"Cataluña"
"Y15-24","ES52",2008,26.2,"Comunidad Valenciana"
"Y15-24","ES53",2008,24.4,"Illes Balears"
"Y15-24","ES6",2008,30,"Sur (ES)"
"Y15-24","ES61",2008,31.1,"Andalucía"
"Y15-24","ES62",2008,23.4,"Región de Murcia"
"Y15-24","ES63",2008,39.6,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2008,38.2,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2008,31.9,"Canarias (ES)"
"Y15-24","ES70",2008,31.9,"Canarias (ES)"
"Y15-24","EU15",2008,15.5,"European Union (15 countries)"
"Y15-24","EU27",2008,15.7,"European Union (27 countries)"
"Y15-24","EU28",2008,15.7,"European Union (28 countries)"
"Y15-24","FI",2008,16.5,"Finland"
"Y15-24","FI1",2008,16.5,"Manner-Suomi"
"Y15-24","FI19",2008,16.1,"Länsi-Suomi"
"Y15-24","FI1B",2008,14.1,"Helsinki-Uusimaa"
"Y15-24","FI1C",2008,15.9,"Etelä-Suomi"
"Y15-24","FI1D",2008,20.4,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2008,NA,"Åland"
"Y15-24","FI20",2008,NA,"Åland"
"Y15-24","FR",2008,19.1,"France"
"Y15-24","FR1",2008,18.6,"Île de France"
"Y15-24","FR10",2008,18.6,"Île de France"
"Y15-24","FR2",2008,18.1,"Bassin Parisien"
"Y15-24","FR21",2008,19.2,"Champagne-Ardenne"
"Y15-24","FR22",2008,17.8,"Picardie"
"Y15-24","FR23",2008,22.1,"Haute-Normandie"
"Y15-24","FR24",2008,14.5,"Centre (FR)"
"Y15-24","FR25",2008,16.4,"Basse-Normandie"
"Y15-24","FR26",2008,18.4,"Bourgogne"
"Y15-24","FR3",2008,27.5,"Nord - Pas-de-Calais"
"Y15-24","FR30",2008,27.5,"Nord - Pas-de-Calais"
"Y15-24","FR4",2008,16.7,"Est (FR)"
"Y15-24","FR41",2008,18.3,"Lorraine"
"Y15-24","FR42",2008,13.8,"Alsace"
"Y15-24","FR43",2008,18.9,"Franche-Comté"
"Y15-24","FR5",2008,16,"Ouest (FR)"
"Y15-24","FR51",2008,16,"Pays de la Loire"
"Y15-24","FR52",2008,14.9,"Bretagne"
"Y15-24","FR53",2008,18.2,"Poitou-Charentes"
"Y15-24","FR6",2008,17.8,"Sud-Ouest (FR)"
"Y15-24","FR61",2008,20.8,"Aquitaine"
"Y15-24","FR62",2008,16.1,"Midi-Pyrénées"
"Y15-24","FR63",2008,NA,"Limousin"
"Y15-24","FR7",2008,13.5,"Centre-Est (FR)"
"Y15-24","FR71",2008,14,"Rhône-Alpes"
"Y15-24","FR72",2008,NA,"Auvergne"
"Y15-24","FR8",2008,22.2,"Méditerranée"
"Y15-24","FR81",2008,26.1,"Languedoc-Roussillon"
"Y15-24","FR82",2008,20.6,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2008,NA,"Corse"
"Y15-24","FR9",2008,48.1,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2008,51.7,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2008,50,"Martinique (NUTS 2010)"
"Y15-24","FR93",2008,39.6,"Guyane (NUTS 2010)"
"Y15-24","FR94",2008,47.6,"Réunion (NUTS 2010)"
"Y15-24","HR",2008,23.7,"Croatia"
"Y15-24","HR0",2008,23.7,"Hrvatska"
"Y15-24","HR03",2008,19.7,"Jadranska Hrvatska"
"Y15-24","HR04",2008,25.4,"Kontinentalna Hrvatska"
"Y15-24","HU",2008,19.5,"Hungary"
"Y15-24","HU1",2008,11.2,"Közép-Magyarország"
"Y15-24","HU10",2008,11.2,"Közép-Magyarország"
"Y15-24","HU2",2008,16.6,"Dunántúl"
"Y15-24","HU21",2008,15.3,"Közép-Dunántúl"
"Y15-24","HU22",2008,10.1,"Nyugat-Dunántúl"
"Y15-24","HU23",2008,25.9,"Dél-Dunántúl"
"Y15-24","HU3",2008,26.5,"Alföld és Észak"
"Y15-24","HU31",2008,29.7,"Észak-Magyarország"
"Y15-24","HU32",2008,28.4,"Észak-Alföld"
"Y15-24","HU33",2008,20.9,"Dél-Alföld"
"Y15-24","IE",2008,13.3,"Ireland"
"Y15-24","IE0",2008,13.3,"Éire/Ireland"
"Y15-24","IE01",2008,15.8,"Border, Midland and Western"
"Y15-24","IE02",2008,12.4,"Southern and Eastern"
"Y15-24","IS",2008,8.2,"Iceland"
"Y15-24","IS0",2008,8.2,"Ísland"
"Y15-24","IS00",2008,8.2,"Ísland"
"Y15-24","IT",2008,21.2,"Italy"
"Y15-24","ITC",2008,13.8,"Nord-Ovest"
"Y15-24","ITC1",2008,15,"Piemonte"
"Y15-24","ITC2",2008,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2008,21.8,"Liguria"
"Y15-24","ITC4",2008,12.3,"Lombardia"
"Y15-24","ITF",2008,31.3,"Sud"
"Y15-24","ITF1",2008,20.5,"Abruzzo"
"Y15-24","ITF2",2008,28.8,"Molise"
"Y15-24","ITF3",2008,32.4,"Campania"
"Y15-24","ITF4",2008,31.6,"Puglia"
"Y15-24","ITF5",2008,34.8,"Basilicata"
"Y15-24","ITF6",2008,34.4,"Calabria"
"Y15-24","ITG",2008,38.5,"Isole"
"Y15-24","ITG1",2008,39.1,"Sicilia"
"Y15-24","ITG2",2008,36.8,"Sardegna"
"Y15-24","ITH",2008,10.5,"Nord-Est"
"Y15-24","ITH1",2008,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2008,8.4,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2008,10.4,"Veneto"
"Y15-24","ITH4",2008,13.2,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2008,11,"Emilia-Romagna"
"Y15-24","ITI",2008,19.5,"Centro (IT)"
"Y15-24","ITI1",2008,14.6,"Toscana"
"Y15-24","ITI2",2008,14.4,"Umbria"
"Y15-24","ITI3",2008,12.5,"Marche"
"Y15-24","ITI4",2008,26.1,"Lazio"
"Y15-24","LT",2008,13.3,"Lithuania"
"Y15-24","LT0",2008,13.3,"Lietuva"
"Y15-24","LT00",2008,13.3,"Lietuva"
"Y15-24","LU",2008,17.9,"Luxembourg"
"Y15-24","LU0",2008,17.9,"Luxembourg"
"Y15-24","LU00",2008,17.9,"Luxembourg"
"Y15-24","LV",2008,13.6,"Latvia"
"Y15-24","LV0",2008,13.6,"Latvija"
"Y15-24","LV00",2008,13.6,"Latvija"
"Y15-24","MK",2008,56.4,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2008,56.4,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2008,56.4,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2008,11.7,"Malta"
"Y15-24","MT0",2008,11.7,"Malta"
"Y15-24","MT00",2008,11.7,"Malta"
"Y15-24","NL",2008,5.3,"Netherlands"
"Y15-24","NL1",2008,6.7,"Noord-Nederland"
"Y15-24","NL11",2008,7.3,"Groningen"
"Y15-24","NL12",2008,5.7,"Friesland (NL)"
"Y15-24","NL13",2008,7.1,"Drenthe"
"Y15-24","NL2",2008,5.1,"Oost-Nederland"
"Y15-24","NL21",2008,4.3,"Overijssel"
"Y15-24","NL22",2008,5.1,"Gelderland"
"Y15-24","NL23",2008,6.7,"Flevoland"
"Y15-24","NL3",2008,5.2,"West-Nederland"
"Y15-24","NL31",2008,4.3,"Utrecht"
"Y15-24","NL32",2008,4.7,"Noord-Holland"
"Y15-24","NL33",2008,6,"Zuid-Holland"
"Y15-24","NL34",2008,NA,"Zeeland"
"Y15-24","NL4",2008,5,"Zuid-Nederland"
"Y15-24","NL41",2008,4.3,"Noord-Brabant"
"Y15-24","NL42",2008,6.6,"Limburg (NL)"
"Y15-24","NO",2008,7.5,"Norway"
"Y15-24","NO0",2008,7.5,"Norge"
"Y15-24","NO01",2008,7.7,"Oslo og Akershus"
"Y15-24","NO02",2008,9.3,"Hedmark og Oppland"
"Y15-24","NO03",2008,9,"Sør-Østlandet"
"Y15-24","NO04",2008,4.1,"Agder og Rogaland"
"Y15-24","NO05",2008,6.4,"Vestlandet"
"Y15-24","NO06",2008,10.3,"Trøndelag"
"Y15-24","NO07",2008,7.9,"Nord-Norge"
"Y15-24","PL",2008,17.3,"Poland"
"Y15-24","PL1",2008,15.5,"Region Centralny"
"Y15-24","PL11",2008,16.8,"Lódzkie"
"Y15-24","PL12",2008,14.9,"Mazowieckie"
"Y15-24","PL2",2008,18,"Region Poludniowy"
"Y15-24","PL21",2008,19,"Malopolskie"
"Y15-24","PL22",2008,17.2,"Slaskie"
"Y15-24","PL3",2008,21.1,"Region Wschodni"
"Y15-24","PL31",2008,24.5,"Lubelskie"
"Y15-24","PL32",2008,21.6,"Podkarpackie"
"Y15-24","PL33",2008,20.2,"Swietokrzyskie"
"Y15-24","PL34",2008,15.3,"Podlaskie"
"Y15-24","PL4",2008,15,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2008,12.7,"Wielkopolskie"
"Y15-24","PL42",2008,21.9,"Zachodniopomorskie"
"Y15-24","PL43",2008,15.7,"Lubuskie"
"Y15-24","PL5",2008,19.1,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2008,19.9,"Dolnoslaskie"
"Y15-24","PL52",2008,16.6,"Opolskie"
"Y15-24","PL6",2008,15.3,"Region Pólnocny"
"Y15-24","PL61",2008,19,"Kujawsko-Pomorskie"
"Y15-24","PL62",2008,16,"Warminsko-Mazurskie"
"Y15-24","PL63",2008,11.3,"Pomorskie"
"Y15-24","PT",2008,16.7,"Portugal"
"Y15-24","PT1",2008,16.8,"Continente"
"Y15-24","PT11",2008,16.4,"Norte"
"Y15-24","PT15",2008,NA,"Algarve"
"Y15-24","PT16",2008,12.1,"Centro (PT)"
"Y15-24","PT17",2008,20.7,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2008,20,"Alentejo"
"Y15-24","PT2",2008,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2008,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2008,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2008,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2008,18.6,"Romania"
"Y15-24","RO1",2008,18.3,"Macroregiunea unu"
"Y15-24","RO11",2008,13.5,"Nord-Vest"
"Y15-24","RO12",2008,22.6,"Centru"
"Y15-24","RO2",2008,17.2,"Macroregiunea doi"
"Y15-24","RO21",2008,14,"Nord-Est"
"Y15-24","RO22",2008,21.7,"Sud-Est"
"Y15-24","RO3",2008,18.8,"Macroregiunea trei"
"Y15-24","RO31",2008,19.4,"Sud - Muntenia"
"Y15-24","RO32",2008,17.4,"Bucuresti - Ilfov"
"Y15-24","RO4",2008,21.1,"Macroregiunea patru"
"Y15-24","RO41",2008,21.7,"Sud-Vest Oltenia"
"Y15-24","RO42",2008,20.4,"Vest"
"Y15-24","SE",2008,20.2,"Sweden"
"Y15-24","SE1",2008,20,"Östra Sverige"
"Y15-24","SE11",2008,18.1,"Stockholm"
"Y15-24","SE12",2008,22.1,"Östra Mellansverige"
"Y15-24","SE2",2008,20.2,"Södra Sverige"
"Y15-24","SE21",2008,16.7,"Småland med öarna"
"Y15-24","SE22",2008,22,"Sydsverige"
"Y15-24","SE23",2008,20.5,"Västsverige"
"Y15-24","SE3",2008,20.6,"Norra Sverige"
"Y15-24","SE31",2008,19,"Norra Mellansverige"
"Y15-24","SE32",2008,27.1,"Mellersta Norrland"
"Y15-24","SE33",2008,18.7,"Övre Norrland"
"Y15-24","SI",2008,10.4,"Slovenia"
"Y15-24","SI0",2008,10.4,"Slovenija"
"Y15-24","SI01",2008,12.2,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2008,8.5,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2008,19,"Slovakia"
"Y15-24","SK0",2008,19,"Slovensko"
"Y15-24","SK01",2008,NA,"Bratislavský kraj"
"Y15-24","SK02",2008,12,"Západné Slovensko"
"Y15-24","SK03",2008,25.3,"Stredné Slovensko"
"Y15-24","SK04",2008,26.9,"Východné Slovensko"
"Y15-24","TR",2008,18.5,"Turkey"
"Y15-24","TR1",2008,16.3,"Istanbul"
"Y15-24","TR10",2008,16.3,"Istanbul"
"Y15-24","TR2",2008,17.7,"Bati Marmara"
"Y15-24","TR21",2008,20.2,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2008,15,"Balikesir, Çanakkale"
"Y15-24","TR3",2008,17.9,"Ege"
"Y15-24","TR31",2008,21,"Izmir"
"Y15-24","TR32",2008,17.8,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2008,13.8,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2008,19.6,"Dogu Marmara"
"Y15-24","TR41",2008,18.6,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2008,20.9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2008,21.3,"Bati Anadolu"
"Y15-24","TR51",2008,22.9,"Ankara"
"Y15-24","TR52",2008,19.1,"Konya, Karaman"
"Y15-24","TR6",2008,20.9,"Akdeniz"
"Y15-24","TR61",2008,16.1,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2008,24.7,"Adana, Mersin"
"Y15-24","TR63",2008,20.8,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2008,22.2,"Orta Anadolu"
"Y15-24","TR71",2008,22,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2008,22.3,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2008,13.4,"Bati Karadeniz"
"Y15-24","TR81",2008,16.3,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2008,10.3,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2008,13.3,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2008,13.2,"Dogu Karadeniz"
"Y15-24","TR90",2008,13.2,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2008,10.2,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2008,10.8,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2008,9.6,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2008,24,"Ortadogu Anadolu"
"Y15-24","TRB1",2008,26.7,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2008,21.5,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2008,21.1,"Güneydogu Anadolu"
"Y15-24","TRC1",2008,22,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2008,17.3,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2008,26,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2008,15,"United Kingdom"
"Y15-24","UKC",2008,18.4,"North East (UK)"
"Y15-24","UKC1",2008,17.3,"Tees Valley and Durham"
"Y15-24","UKC2",2008,19.3,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2008,17.5,"North West (UK)"
"Y15-24","UKD1",2008,NA,"Cumbria"
"Y15-24","UKD3",2008,18.6,"Greater Manchester"
"Y15-24","UKD4",2008,14.2,"Lancashire"
"Y15-24","UKD6",2008,15,"Cheshire"
"Y15-24","UKD7",2008,23.1,"Merseyside"
"Y15-24","UKE",2008,15.4,"Yorkshire and The Humber"
"Y15-24","UKE1",2008,11.3,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2008,10.2,"North Yorkshire"
"Y15-24","UKE3",2008,20.3,"South Yorkshire"
"Y15-24","UKE4",2008,16,"West Yorkshire"
"Y15-24","UKF",2008,15.4,"East Midlands (UK)"
"Y15-24","UKF1",2008,14.3,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2008,16.8,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2008,15.1,"Lincolnshire"
"Y15-24","UKG",2008,16.8,"West Midlands (UK)"
"Y15-24","UKG1",2008,13.9,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2008,10.8,"Shropshire and Staffordshire"
"Y15-24","UKG3",2008,21.7,"West Midlands"
"Y15-24","UKH",2008,13.2,"East of England"
"Y15-24","UKH1",2008,12.7,"East Anglia"
"Y15-24","UKH2",2008,12.8,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2008,14.1,"Essex"
"Y15-24","UKI",2008,19.5,"London"
"Y15-24","UKI1",2008,21.3,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2008,18.3,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2008,12.3,"South East (UK)"
"Y15-24","UKJ1",2008,11.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2008,13.3,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2008,8.8,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2008,16.2,"Kent"
"Y15-24","UKK",2008,10.1,"South West (UK)"
"Y15-24","UKK1",2008,8.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2008,12.2,"Dorset and Somerset"
"Y15-24","UKK3",2008,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2008,11.2,"Devon"
"Y15-24","UKL",2008,16,"Wales"
"Y15-24","UKL1",2008,16.9,"West Wales and The Valleys"
"Y15-24","UKL2",2008,14.1,"East Wales"
"Y15-24","UKM",2008,12.9,"Scotland"
"Y15-24","UKM2",2008,14.7,"Eastern Scotland"
"Y15-24","UKM3",2008,14.1,"South Western Scotland"
"Y15-24","UKM5",2008,NA,"North Eastern Scotland"
"Y15-24","UKM6",2008,NA,"Highlands and Islands"
"Y15-24","UKN",2008,11.7,"Northern Ireland (UK)"
"Y15-24","UKN0",2008,11.7,"Northern Ireland (UK)"
"Y20-64","AT",2008,3.8,"Austria"
"Y20-64","AT1",2008,5,"Ostösterreich"
"Y20-64","AT11",2008,3.8,"Burgenland (AT)"
"Y20-64","AT12",2008,3.4,"Niederösterreich"
"Y20-64","AT13",2008,6.7,"Wien"
"Y20-64","AT2",2008,3.4,"Südösterreich"
"Y20-64","AT21",2008,3.4,"Kärnten"
"Y20-64","AT22",2008,3.4,"Steiermark"
"Y20-64","AT3",2008,2.6,"Westösterreich"
"Y20-64","AT31",2008,2.5,"Oberösterreich"
"Y20-64","AT32",2008,2.5,"Salzburg"
"Y20-64","AT33",2008,2.3,"Tirol"
"Y20-64","AT34",2008,3.8,"Vorarlberg"
"Y20-64","BE",2008,6.8,"Belgium"
"Y20-64","BE1",2008,15.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2008,15.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2008,3.8,"Vlaams Gewest"
"Y20-64","BE21",2008,4.5,"Prov. Antwerpen"
"Y20-64","BE22",2008,4.1,"Prov. Limburg (BE)"
"Y20-64","BE23",2008,3.5,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2008,4.1,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2008,2.6,"Prov. West-Vlaanderen"
"Y20-64","BE3",2008,9.7,"Région wallonne"
"Y20-64","BE31",2008,6.3,"Prov. Brabant Wallon"
"Y20-64","BE32",2008,11.2,"Prov. Hainaut"
"Y20-64","BE33",2008,10.3,"Prov. Liège"
"Y20-64","BE34",2008,7.4,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2008,8.5,"Prov. Namur"
"Y20-64","BG",2008,5.4,"Bulgaria"
"Y20-64","BG3",2008,7.2,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2008,6.9,"Severozapaden"
"Y20-64","BG32",2008,8.4,"Severen tsentralen"
"Y20-64","BG33",2008,8.3,"Severoiztochen"
"Y20-64","BG34",2008,5.5,"Yugoiztochen"
"Y20-64","BG4",2008,3.7,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2008,2.8,"Yugozapaden"
"Y20-64","BG42",2008,4.9,"Yuzhen tsentralen"
"Y20-64","CH",2008,3.2,"Switzerland"
"Y20-64","CH0",2008,3.2,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2008,4.2,"Région lémanique"
"Y20-64","CH02",2008,3.1,"Espace Mittelland"
"Y20-64","CH03",2008,2.9,"Nordwestschweiz"
"Y20-64","CH04",2008,3.1,"Zürich"
"Y20-64","CH05",2008,2.6,"Ostschweiz"
"Y20-64","CH06",2008,2.3,"Zentralschweiz"
"Y20-64","CH07",2008,4.7,"Ticino"
"Y20-64","CY",2008,3.7,"Cyprus"
"Y20-64","CY0",2008,3.7,"Kypros"
"Y20-64","CY00",2008,3.7,"Kypros"
"Y20-64","CZ",2008,4.3,"Czech Republic"
"Y20-64","CZ0",2008,4.3,"Ceská republika"
"Y20-64","CZ01",2008,1.9,"Praha"
"Y20-64","CZ02",2008,2.5,"Strední Cechy"
"Y20-64","CZ03",2008,2.9,"Jihozápad"
"Y20-64","CZ04",2008,7.4,"Severozápad"
"Y20-64","CZ05",2008,3.9,"Severovýchod"
"Y20-64","CZ06",2008,4,"Jihovýchod"
"Y20-64","CZ07",2008,4.8,"Strední Morava"
"Y20-64","CZ08",2008,7.1,"Moravskoslezsko"
"Y20-64","DE",2008,7.5,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2008,4.2,"Baden-Württemberg"
"Y20-64","DE11",2008,4.2,"Stuttgart"
"Y20-64","DE12",2008,4.8,"Karlsruhe"
"Y20-64","DE13",2008,3.7,"Freiburg"
"Y20-64","DE14",2008,3.8,"Tübingen"
"Y20-64","DE2",2008,4.2,"Bayern"
"Y20-64","DE21",2008,3.3,"Oberbayern"
"Y20-64","DE22",2008,4.2,"Niederbayern"
"Y20-64","DE23",2008,4.2,"Oberpfalz"
"Y20-64","DE24",2008,6.1,"Oberfranken"
"Y20-64","DE25",2008,5.5,"Mittelfranken"
"Y20-64","DE26",2008,4.3,"Unterfranken"
"Y20-64","DE27",2008,4,"Schwaben"
"Y20-64","DE3",2008,15.2,"Berlin"
"Y20-64","DE30",2008,15.2,"Berlin"
"Y20-64","DE4",2008,11.6,"Brandenburg"
"Y20-64","DE40",2008,11.6,"Brandenburg"
"Y20-64","DE5",2008,9.6,"Bremen"
"Y20-64","DE50",2008,9.6,"Bremen"
"Y20-64","DE6",2008,6.9,"Hamburg"
"Y20-64","DE60",2008,6.9,"Hamburg"
"Y20-64","DE7",2008,6.4,"Hessen"
"Y20-64","DE71",2008,6.1,"Darmstadt"
"Y20-64","DE72",2008,6.3,"Gießen"
"Y20-64","DE73",2008,7.5,"Kassel"
"Y20-64","DE8",2008,15,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2008,15,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2008,7.1,"Niedersachsen"
"Y20-64","DE91",2008,8.6,"Braunschweig"
"Y20-64","DE92",2008,7.6,"Hannover"
"Y20-64","DE93",2008,6.2,"Lüneburg"
"Y20-64","DE94",2008,6.2,"Weser-Ems"
"Y20-64","DEA",2008,7.3,"Nordrhein-Westfalen"
"Y20-64","DEA1",2008,7.3,"Düsseldorf"
"Y20-64","DEA2",2008,6.9,"Köln"
"Y20-64","DEA3",2008,6.4,"Münster"
"Y20-64","DEA4",2008,6.9,"Detmold"
"Y20-64","DEA5",2008,8.5,"Arnsberg"
"Y20-64","DEB",2008,5.4,"Rheinland-Pfalz"
"Y20-64","DEB1",2008,5.6,"Koblenz"
"Y20-64","DEB2",2008,5.1,"Trier"
"Y20-64","DEB3",2008,5.4,"Rheinhessen-Pfalz"
"Y20-64","DEC",2008,6.8,"Saarland"
"Y20-64","DEC0",2008,6.8,"Saarland"
"Y20-64","DED",2008,13.1,"Sachsen"
"Y20-64","DED2",2008,12.4,"Dresden"
"Y20-64","DED4",2008,12.9,"Chemnitz"
"Y20-64","DED5",2008,14.4,"Leipzig"
"Y20-64","DEE",2008,14.6,"Sachsen-Anhalt"
"Y20-64","DEE0",2008,14.6,"Sachsen-Anhalt"
"Y20-64","DEF",2008,6.7,"Schleswig-Holstein"
"Y20-64","DEF0",2008,6.7,"Schleswig-Holstein"
"Y20-64","DEG",2008,10.8,"Thüringen"
"Y20-64","DEG0",2008,10.8,"Thüringen"
"Y20-64","DK",2008,3,"Denmark"
"Y20-64","DK0",2008,3,"Danmark"
"Y20-64","DK01",2008,3.3,"Hovedstaden"
"Y20-64","DK02",2008,2.8,"Sjælland"
"Y20-64","DK03",2008,2.7,"Syddanmark"
"Y20-64","DK04",2008,2.8,"Midtjylland"
"Y20-64","DK05",2008,3.3,"Nordjylland"
"Y20-64","EA17",2008,7.3,"Euro area (17 countries)"
"Y20-64","EA18",2008,7.3,"Euro area (18 countries)"
"Y20-64","EA19",2008,7.3,"Euro area (19 countries)"
"Y20-64","EE",2008,5.2,"Estonia"
"Y20-64","EE0",2008,5.2,"Eesti"
"Y20-64","EE00",2008,5.2,"Eesti"
"Y20-64","EL",2008,7.7,"Greece"
"Y20-64","EL1",2008,8.8,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2008,8.6,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2008,8.4,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2008,12.3,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2008,8.5,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2008,8.7,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2008,9.9,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2008,8.1,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2008,9.6,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2008,8.6,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2008,7.1,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2008,6.6,"Attiki"
"Y20-64","EL30",2008,6.6,"Attiki"
"Y20-64","EL4",2008,6.7,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2008,4.8,"Voreio Aigaio"
"Y20-64","EL42",2008,8.5,"Notio Aigaio"
"Y20-64","EL43",2008,6.3,"Kriti"
"Y20-64","ES",2008,10.6,"Spain"
"Y20-64","ES1",2008,8.1,"Noroeste (ES)"
"Y20-64","ES11",2008,8.3,"Galicia"
"Y20-64","ES12",2008,8.2,"Principado de Asturias"
"Y20-64","ES13",2008,7,"Cantabria"
"Y20-64","ES2",2008,6.5,"Noreste (ES)"
"Y20-64","ES21",2008,6.3,"País Vasco"
"Y20-64","ES22",2008,6.3,"Comunidad Foral de Navarra"
"Y20-64","ES23",2008,7.3,"La Rioja"
"Y20-64","ES24",2008,6.8,"Aragón"
"Y20-64","ES3",2008,8.1,"Comunidad de Madrid"
"Y20-64","ES30",2008,8.1,"Comunidad de Madrid"
"Y20-64","ES4",2008,10.8,"Centro (ES)"
"Y20-64","ES41",2008,9.1,"Castilla y León"
"Y20-64","ES42",2008,11,"Castilla-la Mancha"
"Y20-64","ES43",2008,14.6,"Extremadura"
"Y20-64","ES5",2008,9.5,"Este (ES)"
"Y20-64","ES51",2008,8.3,"Cataluña"
"Y20-64","ES52",2008,11.2,"Comunidad Valenciana"
"Y20-64","ES53",2008,9.5,"Illes Balears"
"Y20-64","ES6",2008,16.1,"Sur (ES)"
"Y20-64","ES61",2008,16.9,"Andalucía"
"Y20-64","ES62",2008,11.8,"Región de Murcia"
"Y20-64","ES63",2008,16.6,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2008,19.3,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2008,16.6,"Canarias (ES)"
"Y20-64","ES70",2008,16.6,"Canarias (ES)"
"Y20-64","EU15",2008,6.8,"European Union (15 countries)"
"Y20-64","EU27",2008,6.7,"European Union (27 countries)"
"Y20-64","EU28",2008,6.7,"European Union (28 countries)"
"Y20-64","FI",2008,5.6,"Finland"
"Y20-64","FI1",2008,5.6,"Manner-Suomi"
"Y20-64","FI19",2008,5.8,"Länsi-Suomi"
"Y20-64","FI1B",2008,3.9,"Helsinki-Uusimaa"
"Y20-64","FI1C",2008,5.5,"Etelä-Suomi"
"Y20-64","FI1D",2008,7.9,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2008,NA,"Åland"
"Y20-64","FI20",2008,NA,"Åland"
"Y20-64","FR",2008,7.1,"France"
"Y20-64","FR1",2008,6.6,"Île de France"
"Y20-64","FR10",2008,6.6,"Île de France"
"Y20-64","FR2",2008,6.4,"Bassin Parisien"
"Y20-64","FR21",2008,7.1,"Champagne-Ardenne"
"Y20-64","FR22",2008,6.8,"Picardie"
"Y20-64","FR23",2008,7.8,"Haute-Normandie"
"Y20-64","FR24",2008,5.2,"Centre (FR)"
"Y20-64","FR25",2008,6,"Basse-Normandie"
"Y20-64","FR26",2008,6.1,"Bourgogne"
"Y20-64","FR3",2008,10.3,"Nord - Pas-de-Calais"
"Y20-64","FR30",2008,10.3,"Nord - Pas-de-Calais"
"Y20-64","FR4",2008,6.7,"Est (FR)"
"Y20-64","FR41",2008,7.7,"Lorraine"
"Y20-64","FR42",2008,5.6,"Alsace"
"Y20-64","FR43",2008,6.5,"Franche-Comté"
"Y20-64","FR5",2008,5.6,"Ouest (FR)"
"Y20-64","FR51",2008,5.8,"Pays de la Loire"
"Y20-64","FR52",2008,4.8,"Bretagne"
"Y20-64","FR53",2008,6.6,"Poitou-Charentes"
"Y20-64","FR6",2008,6.2,"Sud-Ouest (FR)"
"Y20-64","FR61",2008,6.8,"Aquitaine"
"Y20-64","FR62",2008,5.8,"Midi-Pyrénées"
"Y20-64","FR63",2008,5.1,"Limousin"
"Y20-64","FR7",2008,6.2,"Centre-Est (FR)"
"Y20-64","FR71",2008,6.2,"Rhône-Alpes"
"Y20-64","FR72",2008,6.2,"Auvergne"
"Y20-64","FR8",2008,8,"Méditerranée"
"Y20-64","FR81",2008,9.1,"Languedoc-Roussillon"
"Y20-64","FR82",2008,7.5,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2008,NA,"Corse"
"Y20-64","FR9",2008,22.2,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2008,21.6,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2008,21.7,"Martinique (NUTS 2010)"
"Y20-64","FR93",2008,21,"Guyane (NUTS 2010)"
"Y20-64","FR94",2008,23.1,"Réunion (NUTS 2010)"
"Y20-64","HR",2008,8.1,"Croatia"
"Y20-64","HR0",2008,8.1,"Hrvatska"
"Y20-64","HR03",2008,8.1,"Jadranska Hrvatska"
"Y20-64","HR04",2008,8,"Kontinentalna Hrvatska"
"Y20-64","HU",2008,7.7,"Hungary"
"Y20-64","HU1",2008,4.5,"Közép-Magyarország"
"Y20-64","HU10",2008,4.5,"Közép-Magyarország"
"Y20-64","HU2",2008,6.6,"Dunántúl"
"Y20-64","HU21",2008,5.6,"Közép-Dunántúl"
"Y20-64","HU22",2008,4.9,"Nyugat-Dunántúl"
"Y20-64","HU23",2008,10,"Dél-Dunántúl"
"Y20-64","HU3",2008,11.1,"Alföld és Észak"
"Y20-64","HU31",2008,13.1,"Észak-Magyarország"
"Y20-64","HU32",2008,11.9,"Észak-Alföld"
"Y20-64","HU33",2008,8.6,"Dél-Alföld"
"Y20-64","IE",2008,6.1,"Ireland"
"Y20-64","IE0",2008,6.1,"Éire/Ireland"
"Y20-64","IE01",2008,7,"Border, Midland and Western"
"Y20-64","IE02",2008,5.8,"Southern and Eastern"
"Y20-64","IS",2008,2.2,"Iceland"
"Y20-64","IS0",2008,2.2,"Ísland"
"Y20-64","IS00",2008,2.2,"Ísland"
"Y20-64","IT",2008,6.4,"Italy"
"Y20-64","ITC",2008,4,"Nord-Ovest"
"Y20-64","ITC1",2008,4.9,"Piemonte"
"Y20-64","ITC2",2008,3,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2008,5.1,"Liguria"
"Y20-64","ITC4",2008,3.4,"Lombardia"
"Y20-64","ITF",2008,11,"Sud"
"Y20-64","ITF1",2008,6.6,"Abruzzo"
"Y20-64","ITF2",2008,8.8,"Molise"
"Y20-64","ITF3",2008,12.1,"Campania"
"Y20-64","ITF4",2008,11.1,"Puglia"
"Y20-64","ITF5",2008,10.8,"Basilicata"
"Y20-64","ITF6",2008,11.6,"Calabria"
"Y20-64","ITG",2008,12.7,"Isole"
"Y20-64","ITG1",2008,13.1,"Sicilia"
"Y20-64","ITG2",2008,11.8,"Sardegna"
"Y20-64","ITH",2008,3.2,"Nord-Est"
"Y20-64","ITH1",2008,2.3,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2008,3.1,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2008,3.3,"Veneto"
"Y20-64","ITH4",2008,3.9,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2008,3,"Emilia-Romagna"
"Y20-64","ITI",2008,5.9,"Centro (IT)"
"Y20-64","ITI1",2008,4.9,"Toscana"
"Y20-64","ITI2",2008,4.6,"Umbria"
"Y20-64","ITI3",2008,4.5,"Marche"
"Y20-64","ITI4",2008,7.1,"Lazio"
"Y20-64","LT",2008,5.7,"Lithuania"
"Y20-64","LT0",2008,5.7,"Lietuva"
"Y20-64","LT00",2008,5.7,"Lietuva"
"Y20-64","LU",2008,4.9,"Luxembourg"
"Y20-64","LU0",2008,4.9,"Luxembourg"
"Y20-64","LU00",2008,4.9,"Luxembourg"
"Y20-64","LV",2008,7.6,"Latvia"
"Y20-64","LV0",2008,7.6,"Latvija"
"Y20-64","LV00",2008,7.6,"Latvija"
"Y20-64","MK",2008,33.3,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2008,33.3,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2008,33.3,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2008,4.9,"Malta"
"Y20-64","MT0",2008,4.9,"Malta"
"Y20-64","MT00",2008,4.9,"Malta"
"Y20-64","NL",2008,2.4,"Netherlands"
"Y20-64","NL1",2008,3.1,"Noord-Nederland"
"Y20-64","NL11",2008,3.7,"Groningen"
"Y20-64","NL12",2008,2.4,"Friesland (NL)"
"Y20-64","NL13",2008,3.2,"Drenthe"
"Y20-64","NL2",2008,2.3,"Oost-Nederland"
"Y20-64","NL21",2008,2.2,"Overijssel"
"Y20-64","NL22",2008,2.2,"Gelderland"
"Y20-64","NL23",2008,3,"Flevoland"
"Y20-64","NL3",2008,2.3,"West-Nederland"
"Y20-64","NL31",2008,1.8,"Utrecht"
"Y20-64","NL32",2008,2.2,"Noord-Holland"
"Y20-64","NL33",2008,2.5,"Zuid-Holland"
"Y20-64","NL34",2008,2.4,"Zeeland"
"Y20-64","NL4",2008,2.3,"Zuid-Nederland"
"Y20-64","NL41",2008,2,"Noord-Brabant"
"Y20-64","NL42",2008,2.9,"Limburg (NL)"
"Y20-64","NO",2008,2,"Norway"
"Y20-64","NO0",2008,2,"Norge"
"Y20-64","NO01",2008,2.3,"Oslo og Akershus"
"Y20-64","NO02",2008,1.9,"Hedmark og Oppland"
"Y20-64","NO03",2008,1.9,"Sør-Østlandet"
"Y20-64","NO04",2008,1.5,"Agder og Rogaland"
"Y20-64","NO05",2008,1.6,"Vestlandet"
"Y20-64","NO06",2008,2.6,"Trøndelag"
"Y20-64","NO07",2008,2.3,"Nord-Norge"
"Y20-64","PL",2008,7,"Poland"
"Y20-64","PL1",2008,6.1,"Region Centralny"
"Y20-64","PL11",2008,6.6,"Lódzkie"
"Y20-64","PL12",2008,5.8,"Mazowieckie"
"Y20-64","PL2",2008,6.3,"Region Poludniowy"
"Y20-64","PL21",2008,6.1,"Malopolskie"
"Y20-64","PL22",2008,6.4,"Slaskie"
"Y20-64","PL3",2008,8.4,"Region Wschodni"
"Y20-64","PL31",2008,9,"Lubelskie"
"Y20-64","PL32",2008,8.4,"Podkarpackie"
"Y20-64","PL33",2008,8.8,"Swietokrzyskie"
"Y20-64","PL34",2008,6.5,"Podlaskie"
"Y20-64","PL4",2008,6.9,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2008,6,"Wielkopolskie"
"Y20-64","PL42",2008,9.4,"Zachodniopomorskie"
"Y20-64","PL43",2008,6.3,"Lubuskie"
"Y20-64","PL5",2008,8.4,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2008,9.1,"Dolnoslaskie"
"Y20-64","PL52",2008,6.4,"Opolskie"
"Y20-64","PL6",2008,7.2,"Region Pólnocny"
"Y20-64","PL61",2008,9,"Kujawsko-Pomorskie"
"Y20-64","PL62",2008,7.2,"Warminsko-Mazurskie"
"Y20-64","PL63",2008,5.4,"Pomorskie"
"Y20-64","PT",2008,7.7,"Portugal"
"Y20-64","PT1",2008,7.8,"Continente"
"Y20-64","PT11",2008,8.7,"Norte"
"Y20-64","PT15",2008,7.1,"Algarve"
"Y20-64","PT16",2008,5.9,"Centro (PT)"
"Y20-64","PT17",2008,8.1,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2008,9,"Alentejo"
"Y20-64","PT2",2008,5.2,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2008,5.2,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2008,5.8,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2008,5.8,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2008,5.6,"Romania"
"Y20-64","RO1",2008,5.7,"Macroregiunea unu"
"Y20-64","RO11",2008,3.6,"Nord-Vest"
"Y20-64","RO12",2008,7.9,"Centru"
"Y20-64","RO2",2008,5.6,"Macroregiunea doi"
"Y20-64","RO21",2008,4.6,"Nord-Est"
"Y20-64","RO22",2008,6.9,"Sud-Est"
"Y20-64","RO3",2008,5.2,"Macroregiunea trei"
"Y20-64","RO31",2008,6.6,"Sud - Muntenia"
"Y20-64","RO32",2008,3.2,"Bucuresti - Ilfov"
"Y20-64","RO4",2008,6.1,"Macroregiunea patru"
"Y20-64","RO41",2008,6.7,"Sud-Vest Oltenia"
"Y20-64","RO42",2008,5.4,"Vest"
"Y20-64","SE",2008,5.1,"Sweden"
"Y20-64","SE1",2008,4.8,"Östra Sverige"
"Y20-64","SE11",2008,4.2,"Stockholm"
"Y20-64","SE12",2008,5.7,"Östra Mellansverige"
"Y20-64","SE2",2008,5.1,"Södra Sverige"
"Y20-64","SE21",2008,4.1,"Småland med öarna"
"Y20-64","SE22",2008,6,"Sydsverige"
"Y20-64","SE23",2008,4.8,"Västsverige"
"Y20-64","SE3",2008,5.7,"Norra Sverige"
"Y20-64","SE31",2008,5.7,"Norra Mellansverige"
"Y20-64","SE32",2008,5.5,"Mellersta Norrland"
"Y20-64","SE33",2008,5.7,"Övre Norrland"
"Y20-64","SI",2008,4.3,"Slovenia"
"Y20-64","SI0",2008,4.3,"Slovenija"
"Y20-64","SI01",2008,5.2,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2008,3.3,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2008,9.2,"Slovakia"
"Y20-64","SK0",2008,9.2,"Slovensko"
"Y20-64","SK01",2008,3.3,"Bratislavský kraj"
"Y20-64","SK02",2008,6.3,"Západné Slovensko"
"Y20-64","SK03",2008,12.5,"Stredné Slovensko"
"Y20-64","SK04",2008,12.7,"Východné Slovensko"
"Y20-64","TR",2008,9.4,"Turkey"
"Y20-64","TR1",2008,9.6,"Istanbul"
"Y20-64","TR10",2008,9.6,"Istanbul"
"Y20-64","TR2",2008,7.7,"Bati Marmara"
"Y20-64","TR21",2008,9.5,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2008,5.9,"Balikesir, Çanakkale"
"Y20-64","TR3",2008,9.1,"Ege"
"Y20-64","TR31",2008,10.6,"Izmir"
"Y20-64","TR32",2008,9.4,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2008,6.7,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2008,9.2,"Dogu Marmara"
"Y20-64","TR41",2008,9.3,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2008,9.1,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2008,9.7,"Bati Anadolu"
"Y20-64","TR51",2008,10.1,"Ankara"
"Y20-64","TR52",2008,8.7,"Konya, Karaman"
"Y20-64","TR6",2008,12,"Akdeniz"
"Y20-64","TR61",2008,8.2,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2008,13.8,"Adana, Mersin"
"Y20-64","TR63",2008,14.2,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2008,8.7,"Orta Anadolu"
"Y20-64","TR71",2008,7.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2008,9.3,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2008,5.9,"Bati Karadeniz"
"Y20-64","TR81",2008,5.8,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2008,4.8,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2008,6.2,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2008,4.3,"Dogu Karadeniz"
"Y20-64","TR90",2008,4.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2008,5,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2008,5.3,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2008,4.7,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2008,11.9,"Ortadogu Anadolu"
"Y20-64","TRB1",2008,11.9,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2008,12,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2008,13.7,"Güneydogu Anadolu"
"Y20-64","TRC1",2008,14.5,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2008,12.3,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2008,14.8,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2008,4.8,"United Kingdom"
"Y20-64","UKC",2008,6.2,"North East (UK)"
"Y20-64","UKC1",2008,6.6,"Tees Valley and Durham"
"Y20-64","UKC2",2008,5.9,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2008,5.6,"North West (UK)"
"Y20-64","UKD1",2008,2.7,"Cumbria"
"Y20-64","UKD3",2008,6.4,"Greater Manchester"
"Y20-64","UKD4",2008,4.5,"Lancashire"
"Y20-64","UKD6",2008,4.1,"Cheshire"
"Y20-64","UKD7",2008,7.3,"Merseyside"
"Y20-64","UKE",2008,5,"Yorkshire and The Humber"
"Y20-64","UKE1",2008,4.1,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2008,2.2,"North Yorkshire"
"Y20-64","UKE3",2008,7.1,"South Yorkshire"
"Y20-64","UKE4",2008,5.1,"West Yorkshire"
"Y20-64","UKF",2008,4.7,"East Midlands (UK)"
"Y20-64","UKF1",2008,4.6,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2008,4.8,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2008,4.9,"Lincolnshire"
"Y20-64","UKG",2008,5.6,"West Midlands (UK)"
"Y20-64","UKG1",2008,3.5,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2008,3.6,"Shropshire and Staffordshire"
"Y20-64","UKG3",2008,8.1,"West Midlands"
"Y20-64","UKH",2008,4,"East of England"
"Y20-64","UKH1",2008,3.7,"East Anglia"
"Y20-64","UKH2",2008,4,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2008,4.3,"Essex"
"Y20-64","UKI",2008,6.2,"London"
"Y20-64","UKI1",2008,6.9,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2008,5.8,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2008,3.6,"South East (UK)"
"Y20-64","UKJ1",2008,3.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2008,3.8,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2008,3.1,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2008,4.5,"Kent"
"Y20-64","UKK",2008,3.4,"South West (UK)"
"Y20-64","UKK1",2008,3.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2008,3.3,"Dorset and Somerset"
"Y20-64","UKK3",2008,5.5,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2008,2.8,"Devon"
"Y20-64","UKL",2008,4.8,"Wales"
"Y20-64","UKL1",2008,4.9,"West Wales and The Valleys"
"Y20-64","UKL2",2008,4.7,"East Wales"
"Y20-64","UKM",2008,3.9,"Scotland"
"Y20-64","UKM2",2008,3.9,"Eastern Scotland"
"Y20-64","UKM3",2008,4.7,"South Western Scotland"
"Y20-64","UKM5",2008,2.7,"North Eastern Scotland"
"Y20-64","UKM6",2008,NA,"Highlands and Islands"
"Y20-64","UKN",2008,4,"Northern Ireland (UK)"
"Y20-64","UKN0",2008,4,"Northern Ireland (UK)"
"Y_GE15","AT",2008,4.1,"Austria"
"Y_GE15","AT1",2008,5.4,"Ostösterreich"
"Y_GE15","AT11",2008,4.2,"Burgenland (AT)"
"Y_GE15","AT12",2008,3.7,"Niederösterreich"
"Y_GE15","AT13",2008,7.3,"Wien"
"Y_GE15","AT2",2008,3.7,"Südösterreich"
"Y_GE15","AT21",2008,3.6,"Kärnten"
"Y_GE15","AT22",2008,3.8,"Steiermark"
"Y_GE15","AT3",2008,2.9,"Westösterreich"
"Y_GE15","AT31",2008,2.7,"Oberösterreich"
"Y_GE15","AT32",2008,2.8,"Salzburg"
"Y_GE15","AT33",2008,2.6,"Tirol"
"Y_GE15","AT34",2008,4.1,"Vorarlberg"
"Y_GE15","BE",2008,7,"Belgium"
"Y_GE15","BE1",2008,15.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2008,15.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2008,3.9,"Vlaams Gewest"
"Y_GE15","BE21",2008,4.6,"Prov. Antwerpen"
"Y_GE15","BE22",2008,4.4,"Prov. Limburg (BE)"
"Y_GE15","BE23",2008,3.6,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2008,4.2,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2008,2.7,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2008,10,"Région wallonne"
"Y_GE15","BE31",2008,6.5,"Prov. Brabant Wallon"
"Y_GE15","BE32",2008,11.6,"Prov. Hainaut"
"Y_GE15","BE33",2008,10.5,"Prov. Liège"
"Y_GE15","BE34",2008,7.7,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2008,8.8,"Prov. Namur"
"Y_GE15","BG",2008,5.6,"Bulgaria"
"Y_GE15","BG3",2008,7.5,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2008,7.1,"Severozapaden"
"Y_GE15","BG32",2008,8.5,"Severen tsentralen"
"Y_GE15","BG33",2008,8.6,"Severoiztochen"
"Y_GE15","BG34",2008,5.8,"Yugoiztochen"
"Y_GE15","BG4",2008,3.8,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2008,2.9,"Yugozapaden"
"Y_GE15","BG42",2008,5.1,"Yuzhen tsentralen"
"Y_GE15","CH",2008,3.3,"Switzerland"
"Y_GE15","CH0",2008,3.3,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2008,4.6,"Région lémanique"
"Y_GE15","CH02",2008,3.3,"Espace Mittelland"
"Y_GE15","CH03",2008,3.1,"Nordwestschweiz"
"Y_GE15","CH04",2008,3.1,"Zürich"
"Y_GE15","CH05",2008,2.7,"Ostschweiz"
"Y_GE15","CH06",2008,2.3,"Zentralschweiz"
"Y_GE15","CH07",2008,5,"Ticino"
"Y_GE15","CY",2008,3.7,"Cyprus"
"Y_GE15","CY0",2008,3.7,"Kypros"
"Y_GE15","CY00",2008,3.7,"Kypros"
"Y_GE15","CZ",2008,4.4,"Czech Republic"
"Y_GE15","CZ0",2008,4.4,"Ceská republika"
"Y_GE15","CZ01",2008,1.9,"Praha"
"Y_GE15","CZ02",2008,2.6,"Strední Cechy"
"Y_GE15","CZ03",2008,3.1,"Jihozápad"
"Y_GE15","CZ04",2008,7.8,"Severozápad"
"Y_GE15","CZ05",2008,4,"Severovýchod"
"Y_GE15","CZ06",2008,4,"Jihovýchod"
"Y_GE15","CZ07",2008,4.9,"Strední Morava"
"Y_GE15","CZ08",2008,7.4,"Moravskoslezsko"
"Y_GE15","DE",2008,7.5,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2008,4.2,"Baden-Württemberg"
"Y_GE15","DE11",2008,4.3,"Stuttgart"
"Y_GE15","DE12",2008,4.8,"Karlsruhe"
"Y_GE15","DE13",2008,3.8,"Freiburg"
"Y_GE15","DE14",2008,3.8,"Tübingen"
"Y_GE15","DE2",2008,4.3,"Bayern"
"Y_GE15","DE21",2008,3.4,"Oberbayern"
"Y_GE15","DE22",2008,4.2,"Niederbayern"
"Y_GE15","DE23",2008,4.2,"Oberpfalz"
"Y_GE15","DE24",2008,6.2,"Oberfranken"
"Y_GE15","DE25",2008,5.5,"Mittelfranken"
"Y_GE15","DE26",2008,4.4,"Unterfranken"
"Y_GE15","DE27",2008,4.1,"Schwaben"
"Y_GE15","DE3",2008,15.2,"Berlin"
"Y_GE15","DE30",2008,15.2,"Berlin"
"Y_GE15","DE4",2008,11.5,"Brandenburg"
"Y_GE15","DE40",2008,11.5,"Brandenburg"
"Y_GE15","DE5",2008,9.6,"Bremen"
"Y_GE15","DE50",2008,9.6,"Bremen"
"Y_GE15","DE6",2008,7.1,"Hamburg"
"Y_GE15","DE60",2008,7.1,"Hamburg"
"Y_GE15","DE7",2008,6.5,"Hessen"
"Y_GE15","DE71",2008,6.1,"Darmstadt"
"Y_GE15","DE72",2008,6.6,"Gießen"
"Y_GE15","DE73",2008,7.5,"Kassel"
"Y_GE15","DE8",2008,14.7,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2008,14.7,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2008,7.1,"Niedersachsen"
"Y_GE15","DE91",2008,8.7,"Braunschweig"
"Y_GE15","DE92",2008,7.6,"Hannover"
"Y_GE15","DE93",2008,6.3,"Lüneburg"
"Y_GE15","DE94",2008,6.2,"Weser-Ems"
"Y_GE15","DEA",2008,7.4,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2008,7.4,"Düsseldorf"
"Y_GE15","DEA2",2008,7,"Köln"
"Y_GE15","DEA3",2008,6.4,"Münster"
"Y_GE15","DEA4",2008,7.2,"Detmold"
"Y_GE15","DEA5",2008,8.7,"Arnsberg"
"Y_GE15","DEB",2008,5.6,"Rheinland-Pfalz"
"Y_GE15","DEB1",2008,5.8,"Koblenz"
"Y_GE15","DEB2",2008,5.2,"Trier"
"Y_GE15","DEB3",2008,5.7,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2008,7.1,"Saarland"
"Y_GE15","DEC0",2008,7.1,"Saarland"
"Y_GE15","DED",2008,12.9,"Sachsen"
"Y_GE15","DED2",2008,12.3,"Dresden"
"Y_GE15","DED4",2008,12.7,"Chemnitz"
"Y_GE15","DED5",2008,14.3,"Leipzig"
"Y_GE15","DEE",2008,14.5,"Sachsen-Anhalt"
"Y_GE15","DEE0",2008,14.5,"Sachsen-Anhalt"
"Y_GE15","DEF",2008,6.8,"Schleswig-Holstein"
"Y_GE15","DEF0",2008,6.8,"Schleswig-Holstein"
"Y_GE15","DEG",2008,10.7,"Thüringen"
"Y_GE15","DEG0",2008,10.7,"Thüringen"
"Y_GE15","DK",2008,3.4,"Denmark"
"Y_GE15","DK0",2008,3.4,"Danmark"
"Y_GE15","DK01",2008,3.7,"Hovedstaden"
"Y_GE15","DK02",2008,3.4,"Sjælland"
"Y_GE15","DK03",2008,3.3,"Syddanmark"
"Y_GE15","DK04",2008,3.2,"Midtjylland"
"Y_GE15","DK05",2008,3.7,"Nordjylland"
"Y_GE15","EA17",2008,7.5,"Euro area (17 countries)"
"Y_GE15","EA18",2008,7.5,"Euro area (18 countries)"
"Y_GE15","EA19",2008,7.5,"Euro area (19 countries)"
"Y_GE15","EE",2008,5.5,"Estonia"
"Y_GE15","EE0",2008,5.5,"Eesti"
"Y_GE15","EE00",2008,5.5,"Eesti"
"Y_GE15","EL",2008,7.8,"Greece"
"Y_GE15","EL1",2008,8.8,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2008,8.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2008,8.4,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2008,12.5,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2008,8.3,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2008,8.7,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2008,9.9,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2008,8.3,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2008,9.9,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2008,8.5,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2008,7,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2008,6.7,"Attiki"
"Y_GE15","EL30",2008,6.7,"Attiki"
"Y_GE15","EL4",2008,6.7,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2008,4.7,"Voreio Aigaio"
"Y_GE15","EL42",2008,8.3,"Notio Aigaio"
"Y_GE15","EL43",2008,6.4,"Kriti"
"Y_GE15","ES",2008,11.3,"Spain"
"Y_GE15","ES1",2008,8.4,"Noroeste (ES)"
"Y_GE15","ES11",2008,8.6,"Galicia"
"Y_GE15","ES12",2008,8.5,"Principado de Asturias"
"Y_GE15","ES13",2008,7.2,"Cantabria"
"Y_GE15","ES2",2008,6.9,"Noreste (ES)"
"Y_GE15","ES21",2008,6.6,"País Vasco"
"Y_GE15","ES22",2008,6.8,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2008,7.9,"La Rioja"
"Y_GE15","ES24",2008,7.3,"Aragón"
"Y_GE15","ES3",2008,8.6,"Comunidad de Madrid"
"Y_GE15","ES30",2008,8.6,"Comunidad de Madrid"
"Y_GE15","ES4",2008,11.4,"Centro (ES)"
"Y_GE15","ES41",2008,9.6,"Castilla y León"
"Y_GE15","ES42",2008,11.7,"Castilla-la Mancha"
"Y_GE15","ES43",2008,15.4,"Extremadura"
"Y_GE15","ES5",2008,10.1,"Este (ES)"
"Y_GE15","ES51",2008,8.9,"Cataluña"
"Y_GE15","ES52",2008,12,"Comunidad Valenciana"
"Y_GE15","ES53",2008,10.2,"Illes Balears"
"Y_GE15","ES6",2008,16.9,"Sur (ES)"
"Y_GE15","ES61",2008,17.7,"Andalucía"
"Y_GE15","ES62",2008,12.4,"Región de Murcia"
"Y_GE15","ES63",2008,17.4,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2008,20,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2008,17.2,"Canarias (ES)"
"Y_GE15","ES70",2008,17.2,"Canarias (ES)"
"Y_GE15","EU15",2008,7.1,"European Union (15 countries)"
"Y_GE15","EU27",2008,7,"European Union (27 countries)"
"Y_GE15","EU28",2008,7,"European Union (28 countries)"
"Y_GE15","FI",2008,6.4,"Finland"
"Y_GE15","FI1",2008,6.4,"Manner-Suomi"
"Y_GE15","FI19",2008,6.5,"Länsi-Suomi"
"Y_GE15","FI1B",2008,4.8,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2008,6.2,"Etelä-Suomi"
"Y_GE15","FI1D",2008,8.7,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2008,NA,"Åland"
"Y_GE15","FI20",2008,NA,"Åland"
"Y_GE15","FR",2008,7.5,"France"
"Y_GE15","FR1",2008,6.9,"Île de France"
"Y_GE15","FR10",2008,6.9,"Île de France"
"Y_GE15","FR2",2008,6.8,"Bassin Parisien"
"Y_GE15","FR21",2008,7.5,"Champagne-Ardenne"
"Y_GE15","FR22",2008,7.2,"Picardie"
"Y_GE15","FR23",2008,8.4,"Haute-Normandie"
"Y_GE15","FR24",2008,5.5,"Centre (FR)"
"Y_GE15","FR25",2008,6.3,"Basse-Normandie"
"Y_GE15","FR26",2008,6.4,"Bourgogne"
"Y_GE15","FR3",2008,11,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2008,11,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2008,7,"Est (FR)"
"Y_GE15","FR41",2008,8.1,"Lorraine"
"Y_GE15","FR42",2008,5.9,"Alsace"
"Y_GE15","FR43",2008,6.9,"Franche-Comté"
"Y_GE15","FR5",2008,6,"Ouest (FR)"
"Y_GE15","FR51",2008,6.1,"Pays de la Loire"
"Y_GE15","FR52",2008,5.2,"Bretagne"
"Y_GE15","FR53",2008,7,"Poitou-Charentes"
"Y_GE15","FR6",2008,6.5,"Sud-Ouest (FR)"
"Y_GE15","FR61",2008,7.1,"Aquitaine"
"Y_GE15","FR62",2008,6.1,"Midi-Pyrénées"
"Y_GE15","FR63",2008,5.4,"Limousin"
"Y_GE15","FR7",2008,6.3,"Centre-Est (FR)"
"Y_GE15","FR71",2008,6.3,"Rhône-Alpes"
"Y_GE15","FR72",2008,6.4,"Auvergne"
"Y_GE15","FR8",2008,8.3,"Méditerranée"
"Y_GE15","FR81",2008,9.4,"Languedoc-Roussillon"
"Y_GE15","FR82",2008,7.8,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2008,7.9,"Corse"
"Y_GE15","FR9",2008,23.1,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2008,21.9,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2008,22.3,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2008,21.4,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2008,24.4,"Réunion (NUTS 2010)"
"Y_GE15","HR",2008,8.5,"Croatia"
"Y_GE15","HR0",2008,8.5,"Hrvatska"
"Y_GE15","HR03",2008,8.7,"Jadranska Hrvatska"
"Y_GE15","HR04",2008,8.5,"Kontinentalna Hrvatska"
"Y_GE15","HU",2008,7.8,"Hungary"
"Y_GE15","HU1",2008,4.5,"Közép-Magyarország"
"Y_GE15","HU10",2008,4.5,"Közép-Magyarország"
"Y_GE15","HU2",2008,6.8,"Dunántúl"
"Y_GE15","HU21",2008,5.8,"Közép-Dunántúl"
"Y_GE15","HU22",2008,5,"Nyugat-Dunántúl"
"Y_GE15","HU23",2008,10.3,"Dél-Dunántúl"
"Y_GE15","HU3",2008,11.3,"Alföld és Észak"
"Y_GE15","HU31",2008,13.3,"Észak-Magyarország"
"Y_GE15","HU32",2008,12.1,"Észak-Alföld"
"Y_GE15","HU33",2008,8.7,"Dél-Alföld"
"Y_GE15","IE",2008,6.4,"Ireland"
"Y_GE15","IE0",2008,6.4,"Éire/Ireland"
"Y_GE15","IE01",2008,7.4,"Border, Midland and Western"
"Y_GE15","IE02",2008,6.1,"Southern and Eastern"
"Y_GE15","IS",2008,2.9,"Iceland"
"Y_GE15","IS0",2008,2.9,"Ísland"
"Y_GE15","IS00",2008,2.9,"Ísland"
"Y_GE15","IT",2008,6.7,"Italy"
"Y_GE15","ITC",2008,4.2,"Nord-Ovest"
"Y_GE15","ITC1",2008,5.1,"Piemonte"
"Y_GE15","ITC2",2008,3.3,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2008,5.4,"Liguria"
"Y_GE15","ITC4",2008,3.7,"Lombardia"
"Y_GE15","ITF",2008,11.4,"Sud"
"Y_GE15","ITF1",2008,6.6,"Abruzzo"
"Y_GE15","ITF2",2008,9.1,"Molise"
"Y_GE15","ITF3",2008,12.5,"Campania"
"Y_GE15","ITF4",2008,11.6,"Puglia"
"Y_GE15","ITF5",2008,11,"Basilicata"
"Y_GE15","ITF6",2008,12,"Calabria"
"Y_GE15","ITG",2008,13.3,"Isole"
"Y_GE15","ITG1",2008,13.7,"Sicilia"
"Y_GE15","ITG2",2008,12.2,"Sardegna"
"Y_GE15","ITH",2008,3.4,"Nord-Est"
"Y_GE15","ITH1",2008,2.3,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2008,3.3,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2008,3.4,"Veneto"
"Y_GE15","ITH4",2008,4.3,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2008,3.2,"Emilia-Romagna"
"Y_GE15","ITI",2008,6.1,"Centro (IT)"
"Y_GE15","ITI1",2008,5,"Toscana"
"Y_GE15","ITI2",2008,4.8,"Umbria"
"Y_GE15","ITI3",2008,4.7,"Marche"
"Y_GE15","ITI4",2008,7.5,"Lazio"
"Y_GE15","LT",2008,5.8,"Lithuania"
"Y_GE15","LT0",2008,5.8,"Lietuva"
"Y_GE15","LT00",2008,5.8,"Lietuva"
"Y_GE15","LU",2008,5.1,"Luxembourg"
"Y_GE15","LU0",2008,5.1,"Luxembourg"
"Y_GE15","LU00",2008,5.1,"Luxembourg"
"Y_GE15","LV",2008,7.7,"Latvia"
"Y_GE15","LV0",2008,7.7,"Latvija"
"Y_GE15","LV00",2008,7.7,"Latvija"
"Y_GE15","MK",2008,33.8,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2008,33.8,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2008,33.8,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2008,6,"Malta"
"Y_GE15","MT0",2008,6,"Malta"
"Y_GE15","MT00",2008,6,"Malta"
"Y_GE15","NL",2008,2.8,"Netherlands"
"Y_GE15","NL1",2008,3.4,"Noord-Nederland"
"Y_GE15","NL11",2008,4,"Groningen"
"Y_GE15","NL12",2008,2.9,"Friesland (NL)"
"Y_GE15","NL13",2008,3.6,"Drenthe"
"Y_GE15","NL2",2008,2.7,"Oost-Nederland"
"Y_GE15","NL21",2008,2.6,"Overijssel"
"Y_GE15","NL22",2008,2.6,"Gelderland"
"Y_GE15","NL23",2008,3.4,"Flevoland"
"Y_GE15","NL3",2008,2.7,"West-Nederland"
"Y_GE15","NL31",2008,2.1,"Utrecht"
"Y_GE15","NL32",2008,2.6,"Noord-Holland"
"Y_GE15","NL33",2008,3,"Zuid-Holland"
"Y_GE15","NL34",2008,2.8,"Zeeland"
"Y_GE15","NL4",2008,2.7,"Zuid-Nederland"
"Y_GE15","NL41",2008,2.3,"Noord-Brabant"
"Y_GE15","NL42",2008,3.4,"Limburg (NL)"
"Y_GE15","NO",2008,2.5,"Norway"
"Y_GE15","NO0",2008,2.5,"Norge"
"Y_GE15","NO01",2008,2.9,"Oslo og Akershus"
"Y_GE15","NO02",2008,2.4,"Hedmark og Oppland"
"Y_GE15","NO03",2008,2.7,"Sør-Østlandet"
"Y_GE15","NO04",2008,1.8,"Agder og Rogaland"
"Y_GE15","NO05",2008,2.1,"Vestlandet"
"Y_GE15","NO06",2008,3.3,"Trøndelag"
"Y_GE15","NO07",2008,2.9,"Nord-Norge"
"Y_GE15","PL",2008,7.1,"Poland"
"Y_GE15","PL1",2008,6.2,"Region Centralny"
"Y_GE15","PL11",2008,6.7,"Lódzkie"
"Y_GE15","PL12",2008,6,"Mazowieckie"
"Y_GE15","PL2",2008,6.4,"Region Poludniowy"
"Y_GE15","PL21",2008,6.2,"Malopolskie"
"Y_GE15","PL22",2008,6.6,"Slaskie"
"Y_GE15","PL3",2008,8.2,"Region Wschodni"
"Y_GE15","PL31",2008,8.8,"Lubelskie"
"Y_GE15","PL32",2008,8.2,"Podkarpackie"
"Y_GE15","PL33",2008,8.8,"Swietokrzyskie"
"Y_GE15","PL34",2008,6.4,"Podlaskie"
"Y_GE15","PL4",2008,7,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2008,6.1,"Wielkopolskie"
"Y_GE15","PL42",2008,9.5,"Zachodniopomorskie"
"Y_GE15","PL43",2008,6.5,"Lubuskie"
"Y_GE15","PL5",2008,8.5,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2008,9.1,"Dolnoslaskie"
"Y_GE15","PL52",2008,6.5,"Opolskie"
"Y_GE15","PL6",2008,7.3,"Region Pólnocny"
"Y_GE15","PL61",2008,9.1,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2008,7.4,"Warminsko-Mazurskie"
"Y_GE15","PL63",2008,5.5,"Pomorskie"
"Y_GE15","PT",2008,7.6,"Portugal"
"Y_GE15","PT1",2008,7.6,"Continente"
"Y_GE15","PT11",2008,8.6,"Norte"
"Y_GE15","PT15",2008,7,"Algarve"
"Y_GE15","PT16",2008,5.3,"Centro (PT)"
"Y_GE15","PT17",2008,8.2,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2008,8.9,"Alentejo"
"Y_GE15","PT2",2008,5.4,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2008,5.4,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2008,5.9,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2008,5.9,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2008,5.8,"Romania"
"Y_GE15","RO1",2008,6.1,"Macroregiunea unu"
"Y_GE15","RO11",2008,3.8,"Nord-Vest"
"Y_GE15","RO12",2008,8.5,"Centru"
"Y_GE15","RO2",2008,5.6,"Macroregiunea doi"
"Y_GE15","RO21",2008,4.5,"Nord-Est"
"Y_GE15","RO22",2008,7.2,"Sud-Est"
"Y_GE15","RO3",2008,5.4,"Macroregiunea trei"
"Y_GE15","RO31",2008,6.8,"Sud - Muntenia"
"Y_GE15","RO32",2008,3.4,"Bucuresti - Ilfov"
"Y_GE15","RO4",2008,6.1,"Macroregiunea patru"
"Y_GE15","RO41",2008,6.5,"Sud-Vest Oltenia"
"Y_GE15","RO42",2008,5.7,"Vest"
"Y_GE15","SE",2008,6.2,"Sweden"
"Y_GE15","SE1",2008,5.9,"Östra Sverige"
"Y_GE15","SE11",2008,5.2,"Stockholm"
"Y_GE15","SE12",2008,6.9,"Östra Mellansverige"
"Y_GE15","SE2",2008,6.3,"Södra Sverige"
"Y_GE15","SE21",2008,5,"Småland med öarna"
"Y_GE15","SE22",2008,7.4,"Sydsverige"
"Y_GE15","SE23",2008,6.1,"Västsverige"
"Y_GE15","SE3",2008,6.7,"Norra Sverige"
"Y_GE15","SE31",2008,6.6,"Norra Mellansverige"
"Y_GE15","SE32",2008,7.1,"Mellersta Norrland"
"Y_GE15","SE33",2008,6.6,"Övre Norrland"
"Y_GE15","SI",2008,4.4,"Slovenia"
"Y_GE15","SI0",2008,4.4,"Slovenija"
"Y_GE15","SI01",2008,5.2,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2008,3.4,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2008,9.5,"Slovakia"
"Y_GE15","SK0",2008,9.5,"Slovensko"
"Y_GE15","SK01",2008,3.4,"Bratislavský kraj"
"Y_GE15","SK02",2008,6.4,"Západné Slovensko"
"Y_GE15","SK03",2008,13.1,"Stredné Slovensko"
"Y_GE15","SK04",2008,13.2,"Východné Slovensko"
"Y_GE15","TR",2008,9.7,"Turkey"
"Y_GE15","TR1",2008,10,"Istanbul"
"Y_GE15","TR10",2008,10,"Istanbul"
"Y_GE15","TR2",2008,8.1,"Bati Marmara"
"Y_GE15","TR21",2008,9.9,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2008,6.2,"Balikesir, Çanakkale"
"Y_GE15","TR3",2008,9.4,"Ege"
"Y_GE15","TR31",2008,10.9,"Izmir"
"Y_GE15","TR32",2008,9.6,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2008,7,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2008,9.7,"Dogu Marmara"
"Y_GE15","TR41",2008,9.7,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2008,9.7,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2008,10.2,"Bati Anadolu"
"Y_GE15","TR51",2008,10.8,"Ankara"
"Y_GE15","TR52",2008,9.1,"Konya, Karaman"
"Y_GE15","TR6",2008,12.3,"Akdeniz"
"Y_GE15","TR61",2008,8.5,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2008,14.4,"Adana, Mersin"
"Y_GE15","TR63",2008,14.1,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2008,9.3,"Orta Anadolu"
"Y_GE15","TR71",2008,8.1,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2008,10.1,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2008,6,"Bati Karadeniz"
"Y_GE15","TR81",2008,5.9,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2008,4.9,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2008,6.3,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2008,4.3,"Dogu Karadeniz"
"Y_GE15","TR90",2008,4.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2008,5,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2008,5.2,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2008,4.8,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2008,12.5,"Ortadogu Anadolu"
"Y_GE15","TRB1",2008,12.3,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2008,12.6,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2008,14.4,"Güneydogu Anadolu"
"Y_GE15","TRC1",2008,15,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2008,12.8,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2008,15.8,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2008,5.6,"United Kingdom"
"Y_GE15","UKC",2008,7.5,"North East (UK)"
"Y_GE15","UKC1",2008,7.8,"Tees Valley and Durham"
"Y_GE15","UKC2",2008,7.2,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2008,6.6,"North West (UK)"
"Y_GE15","UKD1",2008,3.1,"Cumbria"
"Y_GE15","UKD3",2008,7.6,"Greater Manchester"
"Y_GE15","UKD4",2008,5.4,"Lancashire"
"Y_GE15","UKD6",2008,5,"Cheshire"
"Y_GE15","UKD7",2008,8.5,"Merseyside"
"Y_GE15","UKE",2008,6,"Yorkshire and The Humber"
"Y_GE15","UKE1",2008,5.1,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2008,2.8,"North Yorkshire"
"Y_GE15","UKE3",2008,8.1,"South Yorkshire"
"Y_GE15","UKE4",2008,6.4,"West Yorkshire"
"Y_GE15","UKF",2008,5.7,"East Midlands (UK)"
"Y_GE15","UKF1",2008,5.2,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2008,6,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2008,6.2,"Lincolnshire"
"Y_GE15","UKG",2008,6.6,"West Midlands (UK)"
"Y_GE15","UKG1",2008,4.3,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2008,4.4,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2008,9.3,"West Midlands"
"Y_GE15","UKH",2008,4.7,"East of England"
"Y_GE15","UKH1",2008,4.5,"East Anglia"
"Y_GE15","UKH2",2008,4.7,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2008,5.1,"Essex"
"Y_GE15","UKI",2008,7.2,"London"
"Y_GE15","UKI1",2008,8,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2008,6.6,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2008,4.3,"South East (UK)"
"Y_GE15","UKJ1",2008,4.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2008,4.4,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2008,3.5,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2008,5.3,"Kent"
"Y_GE15","UKK",2008,4,"South West (UK)"
"Y_GE15","UKK1",2008,3.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2008,4.1,"Dorset and Somerset"
"Y_GE15","UKK3",2008,5.7,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2008,3.8,"Devon"
"Y_GE15","UKL",2008,5.9,"Wales"
"Y_GE15","UKL1",2008,6.1,"West Wales and The Valleys"
"Y_GE15","UKL2",2008,5.6,"East Wales"
"Y_GE15","UKM",2008,4.7,"Scotland"
"Y_GE15","UKM2",2008,4.8,"Eastern Scotland"
"Y_GE15","UKM3",2008,5.4,"South Western Scotland"
"Y_GE15","UKM5",2008,3,"North Eastern Scotland"
"Y_GE15","UKM6",2008,2,"Highlands and Islands"
"Y_GE15","UKN",2008,4.4,"Northern Ireland (UK)"
"Y_GE15","UKN0",2008,4.4,"Northern Ireland (UK)"
"Y_GE25","AT",2008,3.4,"Austria"
"Y_GE25","AT1",2008,4.5,"Ostösterreich"
"Y_GE25","AT11",2008,3.4,"Burgenland (AT)"
"Y_GE25","AT12",2008,2.9,"Niederösterreich"
"Y_GE25","AT13",2008,6.2,"Wien"
"Y_GE25","AT2",2008,3.2,"Südösterreich"
"Y_GE25","AT21",2008,3,"Kärnten"
"Y_GE25","AT22",2008,3.2,"Steiermark"
"Y_GE25","AT3",2008,2.3,"Westösterreich"
"Y_GE25","AT31",2008,2.2,"Oberösterreich"
"Y_GE25","AT32",2008,2.1,"Salzburg"
"Y_GE25","AT33",2008,2,"Tirol"
"Y_GE25","AT34",2008,3.5,"Vorarlberg"
"Y_GE25","BE",2008,5.9,"Belgium"
"Y_GE25","BE1",2008,14.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2008,14.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2008,3.3,"Vlaams Gewest"
"Y_GE25","BE21",2008,4,"Prov. Antwerpen"
"Y_GE25","BE22",2008,3.6,"Prov. Limburg (BE)"
"Y_GE25","BE23",2008,2.8,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2008,3.5,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2008,2.2,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2008,8.2,"Région wallonne"
"Y_GE25","BE31",2008,5.3,"Prov. Brabant Wallon"
"Y_GE25","BE32",2008,9.4,"Prov. Hainaut"
"Y_GE25","BE33",2008,8.9,"Prov. Liège"
"Y_GE25","BE34",2008,5.8,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2008,7.2,"Prov. Namur"
"Y_GE25","BG",2008,5,"Bulgaria"
"Y_GE25","BG3",2008,6.5,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2008,6.1,"Severozapaden"
"Y_GE25","BG32",2008,7.6,"Severen tsentralen"
"Y_GE25","BG33",2008,7.7,"Severoiztochen"
"Y_GE25","BG34",2008,4.9,"Yugoiztochen"
"Y_GE25","BG4",2008,3.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2008,2.6,"Yugozapaden"
"Y_GE25","BG42",2008,4.7,"Yuzhen tsentralen"
"Y_GE25","CH",2008,2.8,"Switzerland"
"Y_GE25","CH0",2008,2.8,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2008,3.6,"Région lémanique"
"Y_GE25","CH02",2008,2.7,"Espace Mittelland"
"Y_GE25","CH03",2008,2.3,"Nordwestschweiz"
"Y_GE25","CH04",2008,2.7,"Zürich"
"Y_GE25","CH05",2008,2.3,"Ostschweiz"
"Y_GE25","CH06",2008,2.2,"Zentralschweiz"
"Y_GE25","CH07",2008,4.1,"Ticino"
"Y_GE25","CY",2008,3.1,"Cyprus"
"Y_GE25","CY0",2008,3.1,"Kypros"
"Y_GE25","CY00",2008,3.1,"Kypros"
"Y_GE25","CZ",2008,3.9,"Czech Republic"
"Y_GE25","CZ0",2008,3.9,"Ceská republika"
"Y_GE25","CZ01",2008,1.7,"Praha"
"Y_GE25","CZ02",2008,2.3,"Strední Cechy"
"Y_GE25","CZ03",2008,2.8,"Jihozápad"
"Y_GE25","CZ04",2008,6.7,"Severozápad"
"Y_GE25","CZ05",2008,3.7,"Severovýchod"
"Y_GE25","CZ06",2008,3.7,"Jihovýchod"
"Y_GE25","CZ07",2008,4.4,"Strední Morava"
"Y_GE25","CZ08",2008,6.7,"Moravskoslezsko"
"Y_GE25","DE",2008,7.1,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2008,3.9,"Baden-Württemberg"
"Y_GE25","DE11",2008,3.9,"Stuttgart"
"Y_GE25","DE12",2008,4.6,"Karlsruhe"
"Y_GE25","DE13",2008,3.4,"Freiburg"
"Y_GE25","DE14",2008,3.3,"Tübingen"
"Y_GE25","DE2",2008,4,"Bayern"
"Y_GE25","DE21",2008,3.2,"Oberbayern"
"Y_GE25","DE22",2008,4.1,"Niederbayern"
"Y_GE25","DE23",2008,4,"Oberpfalz"
"Y_GE25","DE24",2008,5.8,"Oberfranken"
"Y_GE25","DE25",2008,5.3,"Mittelfranken"
"Y_GE25","DE26",2008,4.1,"Unterfranken"
"Y_GE25","DE27",2008,3.8,"Schwaben"
"Y_GE25","DE3",2008,14.9,"Berlin"
"Y_GE25","DE30",2008,14.9,"Berlin"
"Y_GE25","DE4",2008,11.1,"Brandenburg"
"Y_GE25","DE40",2008,11.1,"Brandenburg"
"Y_GE25","DE5",2008,9.5,"Bremen"
"Y_GE25","DE50",2008,9.5,"Bremen"
"Y_GE25","DE6",2008,6.5,"Hamburg"
"Y_GE25","DE60",2008,6.5,"Hamburg"
"Y_GE25","DE7",2008,6,"Hessen"
"Y_GE25","DE71",2008,5.7,"Darmstadt"
"Y_GE25","DE72",2008,5.8,"Gießen"
"Y_GE25","DE73",2008,7.1,"Kassel"
"Y_GE25","DE8",2008,14.6,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2008,14.6,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2008,6.7,"Niedersachsen"
"Y_GE25","DE91",2008,8.3,"Braunschweig"
"Y_GE25","DE92",2008,7.2,"Hannover"
"Y_GE25","DE93",2008,5.7,"Lüneburg"
"Y_GE25","DE94",2008,5.8,"Weser-Ems"
"Y_GE25","DEA",2008,6.9,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2008,6.8,"Düsseldorf"
"Y_GE25","DEA2",2008,6.5,"Köln"
"Y_GE25","DEA3",2008,6.1,"Münster"
"Y_GE25","DEA4",2008,6.6,"Detmold"
"Y_GE25","DEA5",2008,8.2,"Arnsberg"
"Y_GE25","DEB",2008,5.1,"Rheinland-Pfalz"
"Y_GE25","DEB1",2008,5.2,"Koblenz"
"Y_GE25","DEB2",2008,4.4,"Trier"
"Y_GE25","DEB3",2008,5.1,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2008,6.3,"Saarland"
"Y_GE25","DEC0",2008,6.3,"Saarland"
"Y_GE25","DED",2008,12.5,"Sachsen"
"Y_GE25","DED2",2008,11.5,"Dresden"
"Y_GE25","DED4",2008,12.7,"Chemnitz"
"Y_GE25","DED5",2008,13.9,"Leipzig"
"Y_GE25","DEE",2008,14,"Sachsen-Anhalt"
"Y_GE25","DEE0",2008,14,"Sachsen-Anhalt"
"Y_GE25","DEF",2008,6.2,"Schleswig-Holstein"
"Y_GE25","DEF0",2008,6.2,"Schleswig-Holstein"
"Y_GE25","DEG",2008,10.6,"Thüringen"
"Y_GE25","DEG0",2008,10.6,"Thüringen"
"Y_GE25","DK",2008,2.6,"Denmark"
"Y_GE25","DK0",2008,2.6,"Danmark"
"Y_GE25","DK01",2008,3,"Hovedstaden"
"Y_GE25","DK02",2008,2.4,"Sjælland"
"Y_GE25","DK03",2008,2.4,"Syddanmark"
"Y_GE25","DK04",2008,2.2,"Midtjylland"
"Y_GE25","DK05",2008,3,"Nordjylland"
"Y_GE25","EA17",2008,6.5,"Euro area (17 countries)"
"Y_GE25","EA18",2008,6.5,"Euro area (18 countries)"
"Y_GE25","EA19",2008,6.5,"Euro area (19 countries)"
"Y_GE25","EE",2008,4.6,"Estonia"
"Y_GE25","EE0",2008,4.6,"Eesti"
"Y_GE25","EE00",2008,4.6,"Eesti"
"Y_GE25","EL",2008,6.6,"Greece"
"Y_GE25","EL1",2008,7.7,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2008,7.7,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2008,7.4,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2008,10.9,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2008,7.2,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2008,7.1,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2008,8.3,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2008,6.8,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2008,7.7,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2008,6.9,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2008,6,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2008,5.7,"Attiki"
"Y_GE25","EL30",2008,5.7,"Attiki"
"Y_GE25","EL4",2008,6,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2008,3.7,"Voreio Aigaio"
"Y_GE25","EL42",2008,7.7,"Notio Aigaio"
"Y_GE25","EL43",2008,5.8,"Kriti"
"Y_GE25","ES",2008,9.7,"Spain"
"Y_GE25","ES1",2008,7.3,"Noroeste (ES)"
"Y_GE25","ES11",2008,7.5,"Galicia"
"Y_GE25","ES12",2008,7.3,"Principado de Asturias"
"Y_GE25","ES13",2008,6.1,"Cantabria"
"Y_GE25","ES2",2008,5.8,"Noreste (ES)"
"Y_GE25","ES21",2008,5.6,"País Vasco"
"Y_GE25","ES22",2008,5.7,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2008,6.5,"La Rioja"
"Y_GE25","ES24",2008,6,"Aragón"
"Y_GE25","ES3",2008,7.3,"Comunidad de Madrid"
"Y_GE25","ES30",2008,7.3,"Comunidad de Madrid"
"Y_GE25","ES4",2008,9.9,"Centro (ES)"
"Y_GE25","ES41",2008,8.3,"Castilla y León"
"Y_GE25","ES42",2008,10,"Castilla-la Mancha"
"Y_GE25","ES43",2008,13.4,"Extremadura"
"Y_GE25","ES5",2008,8.6,"Este (ES)"
"Y_GE25","ES51",2008,7.6,"Cataluña"
"Y_GE25","ES52",2008,10.2,"Comunidad Valenciana"
"Y_GE25","ES53",2008,8.5,"Illes Balears"
"Y_GE25","ES6",2008,15,"Sur (ES)"
"Y_GE25","ES61",2008,15.8,"Andalucía"
"Y_GE25","ES62",2008,10.8,"Región de Murcia"
"Y_GE25","ES63",2008,14.1,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2008,17.8,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2008,15.5,"Canarias (ES)"
"Y_GE25","ES70",2008,15.5,"Canarias (ES)"
"Y_GE25","EU15",2008,6,"European Union (15 countries)"
"Y_GE25","EU27",2008,5.9,"European Union (27 countries)"
"Y_GE25","EU28",2008,5.9,"European Union (28 countries)"
"Y_GE25","FI",2008,4.9,"Finland"
"Y_GE25","FI1",2008,4.9,"Manner-Suomi"
"Y_GE25","FI19",2008,5.1,"Länsi-Suomi"
"Y_GE25","FI1B",2008,3.4,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2008,4.9,"Etelä-Suomi"
"Y_GE25","FI1D",2008,6.9,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2008,NA,"Åland"
"Y_GE25","FI20",2008,NA,"Åland"
"Y_GE25","FR",2008,6.1,"France"
"Y_GE25","FR1",2008,5.7,"Île de France"
"Y_GE25","FR10",2008,5.7,"Île de France"
"Y_GE25","FR2",2008,5.3,"Bassin Parisien"
"Y_GE25","FR21",2008,6.1,"Champagne-Ardenne"
"Y_GE25","FR22",2008,5.7,"Picardie"
"Y_GE25","FR23",2008,6.1,"Haute-Normandie"
"Y_GE25","FR24",2008,4.5,"Centre (FR)"
"Y_GE25","FR25",2008,5,"Basse-Normandie"
"Y_GE25","FR26",2008,5.1,"Bourgogne"
"Y_GE25","FR3",2008,8.7,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2008,8.7,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2008,5.8,"Est (FR)"
"Y_GE25","FR41",2008,6.9,"Lorraine"
"Y_GE25","FR42",2008,4.9,"Alsace"
"Y_GE25","FR43",2008,5.4,"Franche-Comté"
"Y_GE25","FR5",2008,4.8,"Ouest (FR)"
"Y_GE25","FR51",2008,4.9,"Pays de la Loire"
"Y_GE25","FR52",2008,4,"Bretagne"
"Y_GE25","FR53",2008,5.8,"Poitou-Charentes"
"Y_GE25","FR6",2008,5.3,"Sud-Ouest (FR)"
"Y_GE25","FR61",2008,5.9,"Aquitaine"
"Y_GE25","FR62",2008,5,"Midi-Pyrénées"
"Y_GE25","FR63",2008,4.5,"Limousin"
"Y_GE25","FR7",2008,5.5,"Centre-Est (FR)"
"Y_GE25","FR71",2008,5.4,"Rhône-Alpes"
"Y_GE25","FR72",2008,5.9,"Auvergne"
"Y_GE25","FR8",2008,6.9,"Méditerranée"
"Y_GE25","FR81",2008,7.7,"Languedoc-Roussillon"
"Y_GE25","FR82",2008,6.4,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2008,NA,"Corse"
"Y_GE25","FR9",2008,19.9,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2008,19.5,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2008,19.4,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2008,19.4,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2008,20.4,"Réunion (NUTS 2010)"
"Y_GE25","HR",2008,6.9,"Croatia"
"Y_GE25","HR0",2008,6.9,"Hrvatska"
"Y_GE25","HR03",2008,7.5,"Jadranska Hrvatska"
"Y_GE25","HR04",2008,6.5,"Kontinentalna Hrvatska"
"Y_GE25","HU",2008,6.9,"Hungary"
"Y_GE25","HU1",2008,4.1,"Közép-Magyarország"
"Y_GE25","HU10",2008,4.1,"Közép-Magyarország"
"Y_GE25","HU2",2008,5.9,"Dunántúl"
"Y_GE25","HU21",2008,5,"Közép-Dunántúl"
"Y_GE25","HU22",2008,4.5,"Nyugat-Dunántúl"
"Y_GE25","HU23",2008,8.9,"Dél-Dunántúl"
"Y_GE25","HU3",2008,10,"Alföld és Észak"
"Y_GE25","HU31",2008,11.9,"Észak-Magyarország"
"Y_GE25","HU32",2008,10.6,"Észak-Alföld"
"Y_GE25","HU33",2008,7.7,"Dél-Alföld"
"Y_GE25","IE",2008,5.1,"Ireland"
"Y_GE25","IE0",2008,5.1,"Éire/Ireland"
"Y_GE25","IE01",2008,5.8,"Border, Midland and Western"
"Y_GE25","IE02",2008,4.9,"Southern and Eastern"
"Y_GE25","IS",2008,1.9,"Iceland"
"Y_GE25","IS0",2008,1.9,"Ísland"
"Y_GE25","IS00",2008,1.9,"Ísland"
"Y_GE25","IT",2008,5.6,"Italy"
"Y_GE25","ITC",2008,3.5,"Nord-Ovest"
"Y_GE25","ITC1",2008,4.4,"Piemonte"
"Y_GE25","ITC2",2008,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2008,4.3,"Liguria"
"Y_GE25","ITC4",2008,3,"Lombardia"
"Y_GE25","ITF",2008,9.4,"Sud"
"Y_GE25","ITF1",2008,5.5,"Abruzzo"
"Y_GE25","ITF2",2008,7.4,"Molise"
"Y_GE25","ITF3",2008,10.5,"Campania"
"Y_GE25","ITF4",2008,9.4,"Puglia"
"Y_GE25","ITF5",2008,9,"Basilicata"
"Y_GE25","ITF6",2008,10,"Calabria"
"Y_GE25","ITG",2008,10.8,"Isole"
"Y_GE25","ITG1",2008,11.2,"Sicilia"
"Y_GE25","ITG2",2008,10,"Sardegna"
"Y_GE25","ITH",2008,2.8,"Nord-Est"
"Y_GE25","ITH1",2008,2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2008,2.8,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2008,2.9,"Veneto"
"Y_GE25","ITH4",2008,3.7,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2008,2.7,"Emilia-Romagna"
"Y_GE25","ITI",2008,5.2,"Centro (IT)"
"Y_GE25","ITI1",2008,4.4,"Toscana"
"Y_GE25","ITI2",2008,4,"Umbria"
"Y_GE25","ITI3",2008,4.1,"Marche"
"Y_GE25","ITI4",2008,6.2,"Lazio"
"Y_GE25","LT",2008,5,"Lithuania"
"Y_GE25","LT0",2008,5,"Lietuva"
"Y_GE25","LT00",2008,5,"Lietuva"
"Y_GE25","LU",2008,4,"Luxembourg"
"Y_GE25","LU0",2008,4,"Luxembourg"
"Y_GE25","LU00",2008,4,"Luxembourg"
"Y_GE25","LV",2008,6.9,"Latvia"
"Y_GE25","LV0",2008,6.9,"Latvija"
"Y_GE25","LV00",2008,6.9,"Latvija"
"Y_GE25","MK",2008,30.5,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2008,30.5,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2008,30.5,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2008,4.8,"Malta"
"Y_GE25","MT0",2008,4.8,"Malta"
"Y_GE25","MT00",2008,4.8,"Malta"
"Y_GE25","NL",2008,2.3,"Netherlands"
"Y_GE25","NL1",2008,2.8,"Noord-Nederland"
"Y_GE25","NL11",2008,3.2,"Groningen"
"Y_GE25","NL12",2008,2.3,"Friesland (NL)"
"Y_GE25","NL13",2008,2.9,"Drenthe"
"Y_GE25","NL2",2008,2.2,"Oost-Nederland"
"Y_GE25","NL21",2008,2.2,"Overijssel"
"Y_GE25","NL22",2008,2.1,"Gelderland"
"Y_GE25","NL23",2008,2.7,"Flevoland"
"Y_GE25","NL3",2008,2.2,"West-Nederland"
"Y_GE25","NL31",2008,1.6,"Utrecht"
"Y_GE25","NL32",2008,2.2,"Noord-Holland"
"Y_GE25","NL33",2008,2.4,"Zuid-Holland"
"Y_GE25","NL34",2008,2.6,"Zeeland"
"Y_GE25","NL4",2008,2.2,"Zuid-Nederland"
"Y_GE25","NL41",2008,1.9,"Noord-Brabant"
"Y_GE25","NL42",2008,2.8,"Limburg (NL)"
"Y_GE25","NO",2008,1.7,"Norway"
"Y_GE25","NO0",2008,1.7,"Norge"
"Y_GE25","NO01",2008,2.2,"Oslo og Akershus"
"Y_GE25","NO02",2008,1.4,"Hedmark og Oppland"
"Y_GE25","NO03",2008,1.6,"Sør-Østlandet"
"Y_GE25","NO04",2008,1.4,"Agder og Rogaland"
"Y_GE25","NO05",2008,1.4,"Vestlandet"
"Y_GE25","NO06",2008,2.1,"Trøndelag"
"Y_GE25","NO07",2008,1.9,"Nord-Norge"
"Y_GE25","PL",2008,5.9,"Poland"
"Y_GE25","PL1",2008,5.2,"Region Centralny"
"Y_GE25","PL11",2008,5.6,"Lódzkie"
"Y_GE25","PL12",2008,4.9,"Mazowieckie"
"Y_GE25","PL2",2008,5,"Region Poludniowy"
"Y_GE25","PL21",2008,4.5,"Malopolskie"
"Y_GE25","PL22",2008,5.4,"Slaskie"
"Y_GE25","PL3",2008,6.7,"Region Wschodni"
"Y_GE25","PL31",2008,7.2,"Lubelskie"
"Y_GE25","PL32",2008,6.7,"Podkarpackie"
"Y_GE25","PL33",2008,7.3,"Swietokrzyskie"
"Y_GE25","PL34",2008,5.2,"Podlaskie"
"Y_GE25","PL4",2008,6.1,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2008,5.2,"Wielkopolskie"
"Y_GE25","PL42",2008,8.4,"Zachodniopomorskie"
"Y_GE25","PL43",2008,5.6,"Lubuskie"
"Y_GE25","PL5",2008,7.2,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2008,7.8,"Dolnoslaskie"
"Y_GE25","PL52",2008,5.3,"Opolskie"
"Y_GE25","PL6",2008,6.3,"Region Pólnocny"
"Y_GE25","PL61",2008,7.9,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2008,6.4,"Warminsko-Mazurskie"
"Y_GE25","PL63",2008,4.8,"Pomorskie"
"Y_GE25","PT",2008,6.7,"Portugal"
"Y_GE25","PT1",2008,6.8,"Continente"
"Y_GE25","PT11",2008,7.7,"Norte"
"Y_GE25","PT15",2008,5.9,"Algarve"
"Y_GE25","PT16",2008,4.8,"Centro (PT)"
"Y_GE25","PT17",2008,7.2,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2008,7.9,"Alentejo"
"Y_GE25","PT2",2008,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2008,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2008,4.9,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2008,4.9,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2008,4.4,"Romania"
"Y_GE25","RO1",2008,4.8,"Macroregiunea unu"
"Y_GE25","RO11",2008,2.9,"Nord-Vest"
"Y_GE25","RO12",2008,6.9,"Centru"
"Y_GE25","RO2",2008,4.3,"Macroregiunea doi"
"Y_GE25","RO21",2008,3.5,"Nord-Est"
"Y_GE25","RO22",2008,5.6,"Sud-Est"
"Y_GE25","RO3",2008,4,"Macroregiunea trei"
"Y_GE25","RO31",2008,5.2,"Sud - Muntenia"
"Y_GE25","RO32",2008,2.3,"Bucuresti - Ilfov"
"Y_GE25","RO4",2008,4.7,"Macroregiunea patru"
"Y_GE25","RO41",2008,5,"Sud-Vest Oltenia"
"Y_GE25","RO42",2008,4.2,"Vest"
"Y_GE25","SE",2008,4.1,"Sweden"
"Y_GE25","SE1",2008,4,"Östra Sverige"
"Y_GE25","SE11",2008,3.6,"Stockholm"
"Y_GE25","SE12",2008,4.5,"Östra Mellansverige"
"Y_GE25","SE2",2008,4.1,"Södra Sverige"
"Y_GE25","SE21",2008,3.1,"Småland med öarna"
"Y_GE25","SE22",2008,5.1,"Sydsverige"
"Y_GE25","SE23",2008,3.8,"Västsverige"
"Y_GE25","SE3",2008,4.6,"Norra Sverige"
"Y_GE25","SE31",2008,4.7,"Norra Mellansverige"
"Y_GE25","SE32",2008,4.2,"Mellersta Norrland"
"Y_GE25","SE33",2008,4.8,"Övre Norrland"
"Y_GE25","SI",2008,3.7,"Slovenia"
"Y_GE25","SI0",2008,3.7,"Slovenija"
"Y_GE25","SI01",2008,4.4,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2008,2.8,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2008,8.4,"Slovakia"
"Y_GE25","SK0",2008,8.4,"Slovensko"
"Y_GE25","SK01",2008,3.1,"Bratislavský kraj"
"Y_GE25","SK02",2008,5.8,"Západné Slovensko"
"Y_GE25","SK03",2008,11.7,"Stredné Slovensko"
"Y_GE25","SK04",2008,11.6,"Východné Slovensko"
"Y_GE25","TR",2008,7.8,"Turkey"
"Y_GE25","TR1",2008,8.5,"Istanbul"
"Y_GE25","TR10",2008,8.5,"Istanbul"
"Y_GE25","TR2",2008,6.3,"Bati Marmara"
"Y_GE25","TR21",2008,7.9,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2008,4.7,"Balikesir, Çanakkale"
"Y_GE25","TR3",2008,7.6,"Ege"
"Y_GE25","TR31",2008,8.9,"Izmir"
"Y_GE25","TR32",2008,7.9,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2008,5.5,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2008,7.5,"Dogu Marmara"
"Y_GE25","TR41",2008,7.6,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2008,7.2,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2008,7.8,"Bati Anadolu"
"Y_GE25","TR51",2008,8.5,"Ankara"
"Y_GE25","TR52",2008,6.5,"Konya, Karaman"
"Y_GE25","TR6",2008,10.4,"Akdeniz"
"Y_GE25","TR61",2008,7,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2008,12,"Adana, Mersin"
"Y_GE25","TR63",2008,12.3,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2008,6.8,"Orta Anadolu"
"Y_GE25","TR71",2008,5.6,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2008,7.5,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2008,4.4,"Bati Karadeniz"
"Y_GE25","TR81",2008,4.1,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2008,3.7,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2008,4.7,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2008,2.8,"Dogu Karadeniz"
"Y_GE25","TR90",2008,2.8,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2008,3.9,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2008,4,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2008,3.8,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2008,9.6,"Ortadogu Anadolu"
"Y_GE25","TRB1",2008,9.2,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2008,10,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2008,12,"Güneydogu Anadolu"
"Y_GE25","TRC1",2008,12.3,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2008,11.3,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2008,12.7,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2008,3.9,"United Kingdom"
"Y_GE25","UKC",2008,5.4,"North East (UK)"
"Y_GE25","UKC1",2008,6,"Tees Valley and Durham"
"Y_GE25","UKC2",2008,4.9,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2008,4.6,"North West (UK)"
"Y_GE25","UKD1",2008,2.1,"Cumbria"
"Y_GE25","UKD3",2008,5.2,"Greater Manchester"
"Y_GE25","UKD4",2008,3.7,"Lancashire"
"Y_GE25","UKD6",2008,3.4,"Cheshire"
"Y_GE25","UKD7",2008,6.1,"Merseyside"
"Y_GE25","UKE",2008,4.1,"Yorkshire and The Humber"
"Y_GE25","UKE1",2008,3.8,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2008,1.6,"North Yorkshire"
"Y_GE25","UKE3",2008,5.7,"South Yorkshire"
"Y_GE25","UKE4",2008,4.3,"West Yorkshire"
"Y_GE25","UKF",2008,3.9,"East Midlands (UK)"
"Y_GE25","UKF1",2008,3.7,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2008,4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2008,4.4,"Lincolnshire"
"Y_GE25","UKG",2008,4.7,"West Midlands (UK)"
"Y_GE25","UKG1",2008,3,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2008,3.1,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2008,6.8,"West Midlands"
"Y_GE25","UKH",2008,3.3,"East of England"
"Y_GE25","UKH1",2008,3.1,"East Anglia"
"Y_GE25","UKH2",2008,3.5,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2008,3.5,"Essex"
"Y_GE25","UKI",2008,5.2,"London"
"Y_GE25","UKI1",2008,5.9,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2008,4.8,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2008,2.9,"South East (UK)"
"Y_GE25","UKJ1",2008,2.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2008,2.9,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2008,2.6,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2008,3.6,"Kent"
"Y_GE25","UKK",2008,2.9,"South West (UK)"
"Y_GE25","UKK1",2008,2.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2008,2.7,"Dorset and Somerset"
"Y_GE25","UKK3",2008,4.9,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2008,2.3,"Devon"
"Y_GE25","UKL",2008,4,"Wales"
"Y_GE25","UKL1",2008,3.8,"West Wales and The Valleys"
"Y_GE25","UKL2",2008,4.2,"East Wales"
"Y_GE25","UKM",2008,3.1,"Scotland"
"Y_GE25","UKM2",2008,3,"Eastern Scotland"
"Y_GE25","UKM3",2008,3.8,"South Western Scotland"
"Y_GE25","UKM5",2008,2.3,"North Eastern Scotland"
"Y_GE25","UKM6",2008,NA,"Highlands and Islands"
"Y_GE25","UKN",2008,3,"Northern Ireland (UK)"
"Y_GE25","UKN0",2008,3,"Northern Ireland (UK)"
"Y15-24","AT",2007,9.4,"Austria"
"Y15-24","AT1",2007,12.2,"Ostösterreich"
"Y15-24","AT11",2007,NA,"Burgenland (AT)"
"Y15-24","AT12",2007,8.4,"Niederösterreich"
"Y15-24","AT13",2007,17,"Wien"
"Y15-24","AT2",2007,8.9,"Südösterreich"
"Y15-24","AT21",2007,8.6,"Kärnten"
"Y15-24","AT22",2007,9,"Steiermark"
"Y15-24","AT3",2007,7,"Westösterreich"
"Y15-24","AT31",2007,6.9,"Oberösterreich"
"Y15-24","AT32",2007,NA,"Salzburg"
"Y15-24","AT33",2007,6.9,"Tirol"
"Y15-24","AT34",2007,NA,"Vorarlberg"
"Y15-24","BE",2007,18.8,"Belgium"
"Y15-24","BE1",2007,34.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2007,34.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2007,11.7,"Vlaams Gewest"
"Y15-24","BE21",2007,10.1,"Prov. Antwerpen"
"Y15-24","BE22",2007,12.6,"Prov. Limburg (BE)"
"Y15-24","BE23",2007,13.8,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2007,14.4,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2007,9,"Prov. West-Vlaanderen"
"Y15-24","BE3",2007,27.8,"Région wallonne"
"Y15-24","BE31",2007,19.8,"Prov. Brabant Wallon"
"Y15-24","BE32",2007,34.5,"Prov. Hainaut"
"Y15-24","BE33",2007,25.7,"Prov. Liège"
"Y15-24","BE34",2007,17.3,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2007,25.2,"Prov. Namur"
"Y15-24","BG",2007,15.1,"Bulgaria"
"Y15-24","BG3",2007,20.6,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2007,22.3,"Severozapaden"
"Y15-24","BG32",2007,21.1,"Severen tsentralen"
"Y15-24","BG33",2007,25,"Severoiztochen"
"Y15-24","BG34",2007,14.5,"Yugoiztochen"
"Y15-24","BG4",2007,9.5,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2007,7.1,"Yugozapaden"
"Y15-24","BG42",2007,13.8,"Yuzhen tsentralen"
"Y15-24","CH",2007,7.1,"Switzerland"
"Y15-24","CH0",2007,7.1,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2007,9.2,"Région lémanique"
"Y15-24","CH02",2007,9.1,"Espace Mittelland"
"Y15-24","CH03",2007,5.7,"Nordwestschweiz"
"Y15-24","CH04",2007,6.9,"Zürich"
"Y15-24","CH05",2007,4.7,"Ostschweiz"
"Y15-24","CH06",2007,4.6,"Zentralschweiz"
"Y15-24","CH07",2007,NA,"Ticino"
"Y15-24","CY",2007,10.2,"Cyprus"
"Y15-24","CY0",2007,10.2,"Kypros"
"Y15-24","CY00",2007,10.2,"Kypros"
"Y15-24","CZ",2007,10.7,"Czech Republic"
"Y15-24","CZ0",2007,10.7,"Ceská republika"
"Y15-24","CZ01",2007,6.6,"Praha"
"Y15-24","CZ02",2007,7.5,"Strední Cechy"
"Y15-24","CZ03",2007,6,"Jihozápad"
"Y15-24","CZ04",2007,19.3,"Severozápad"
"Y15-24","CZ05",2007,9.9,"Severovýchod"
"Y15-24","CZ06",2007,11.3,"Jihovýchod"
"Y15-24","CZ07",2007,8.8,"Strední Morava"
"Y15-24","CZ08",2007,15.2,"Moravskoslezsko"
"Y15-24","DE",2007,11.9,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2007,6.8,"Baden-Württemberg"
"Y15-24","DE11",2007,7.6,"Stuttgart"
"Y15-24","DE12",2007,7.3,"Karlsruhe"
"Y15-24","DE13",2007,5.1,"Freiburg"
"Y15-24","DE14",2007,6.7,"Tübingen"
"Y15-24","DE2",2007,8,"Bayern"
"Y15-24","DE21",2007,6.6,"Oberbayern"
"Y15-24","DE22",2007,7,"Niederbayern"
"Y15-24","DE23",2007,7.5,"Oberpfalz"
"Y15-24","DE24",2007,11.3,"Oberfranken"
"Y15-24","DE25",2007,9.8,"Mittelfranken"
"Y15-24","DE26",2007,10.6,"Unterfranken"
"Y15-24","DE27",2007,6.5,"Schwaben"
"Y15-24","DE3",2007,21.2,"Berlin"
"Y15-24","DE30",2007,21.2,"Berlin"
"Y15-24","DE4",2007,17.1,"Brandenburg"
"Y15-24","DE40",2007,17.1,"Brandenburg"
"Y15-24","DE5",2007,NA,"Bremen"
"Y15-24","DE50",2007,NA,"Bremen"
"Y15-24","DE6",2007,11.6,"Hamburg"
"Y15-24","DE60",2007,11.6,"Hamburg"
"Y15-24","DE7",2007,11.9,"Hessen"
"Y15-24","DE71",2007,11.3,"Darmstadt"
"Y15-24","DE72",2007,12.7,"Gießen"
"Y15-24","DE73",2007,12.9,"Kassel"
"Y15-24","DE8",2007,19.4,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2007,19.4,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2007,12.1,"Niedersachsen"
"Y15-24","DE91",2007,13.5,"Braunschweig"
"Y15-24","DE92",2007,13.9,"Hannover"
"Y15-24","DE93",2007,10.9,"Lüneburg"
"Y15-24","DE94",2007,10.5,"Weser-Ems"
"Y15-24","DEA",2007,12.5,"Nordrhein-Westfalen"
"Y15-24","DEA1",2007,14.6,"Düsseldorf"
"Y15-24","DEA2",2007,11.3,"Köln"
"Y15-24","DEA3",2007,9.2,"Münster"
"Y15-24","DEA4",2007,11.3,"Detmold"
"Y15-24","DEA5",2007,14.5,"Arnsberg"
"Y15-24","DEB",2007,10.4,"Rheinland-Pfalz"
"Y15-24","DEB1",2007,9.3,"Koblenz"
"Y15-24","DEB2",2007,NA,"Trier"
"Y15-24","DEB3",2007,12,"Rheinhessen-Pfalz"
"Y15-24","DEC",2007,NA,"Saarland"
"Y15-24","DEC0",2007,NA,"Saarland"
"Y15-24","DED",2007,15.9,"Sachsen"
"Y15-24","DED2",2007,16,"Dresden"
"Y15-24","DED4",2007,14,"Chemnitz"
"Y15-24","DED5",2007,18.4,"Leipzig"
"Y15-24","DEE",2007,19.2,"Sachsen-Anhalt"
"Y15-24","DEE0",2007,19.2,"Sachsen-Anhalt"
"Y15-24","DEF",2007,12.9,"Schleswig-Holstein"
"Y15-24","DEF0",2007,12.9,"Schleswig-Holstein"
"Y15-24","DEG",2007,15,"Thüringen"
"Y15-24","DEG0",2007,15,"Thüringen"
"Y15-24","DK",2007,7.5,"Denmark"
"Y15-24","DK0",2007,7.5,"Danmark"
"Y15-24","DK01",2007,7.1,"Hovedstaden"
"Y15-24","DK02",2007,8,"Sjælland"
"Y15-24","DK03",2007,8,"Syddanmark"
"Y15-24","DK04",2007,6.7,"Midtjylland"
"Y15-24","DK05",2007,8.8,"Nordjylland"
"Y15-24","EA17",2007,15.2,"Euro area (17 countries)"
"Y15-24","EA18",2007,15.2,"Euro area (18 countries)"
"Y15-24","EA19",2007,15.1,"Euro area (19 countries)"
"Y15-24","EE",2007,10.1,"Estonia"
"Y15-24","EE0",2007,10.1,"Eesti"
"Y15-24","EE00",2007,10.1,"Eesti"
"Y15-24","EL",2007,22.7,"Greece"
"Y15-24","EL1",2007,24.7,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2007,25.4,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2007,24.2,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2007,35.7,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2007,22.6,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2007,28,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2007,30.9,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2007,24,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2007,31.7,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2007,25.6,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2007,25.7,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2007,20,"Attiki"
"Y15-24","EL30",2007,20,"Attiki"
"Y15-24","EL4",2007,16.8,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2007,36.4,"Voreio Aigaio"
"Y15-24","EL42",2007,12.5,"Notio Aigaio"
"Y15-24","EL43",2007,14,"Kriti"
"Y15-24","ES",2007,18.1,"Spain"
"Y15-24","ES1",2007,16.3,"Noroeste (ES)"
"Y15-24","ES11",2007,15.9,"Galicia"
"Y15-24","ES12",2007,18.9,"Principado de Asturias"
"Y15-24","ES13",2007,13.8,"Cantabria"
"Y15-24","ES2",2007,15.2,"Noreste (ES)"
"Y15-24","ES21",2007,17.5,"País Vasco"
"Y15-24","ES22",2007,11.8,"Comunidad Foral de Navarra"
"Y15-24","ES23",2007,16.6,"La Rioja"
"Y15-24","ES24",2007,13.7,"Aragón"
"Y15-24","ES3",2007,16.8,"Comunidad de Madrid"
"Y15-24","ES30",2007,16.8,"Comunidad de Madrid"
"Y15-24","ES4",2007,18.5,"Centro (ES)"
"Y15-24","ES41",2007,17.3,"Castilla y León"
"Y15-24","ES42",2007,15.8,"Castilla-la Mancha"
"Y15-24","ES43",2007,26.2,"Extremadura"
"Y15-24","ES5",2007,15.7,"Este (ES)"
"Y15-24","ES51",2007,13.4,"Cataluña"
"Y15-24","ES52",2007,19.1,"Comunidad Valenciana"
"Y15-24","ES53",2007,15.2,"Illes Balears"
"Y15-24","ES6",2007,22.4,"Sur (ES)"
"Y15-24","ES61",2007,23.2,"Andalucía"
"Y15-24","ES62",2007,16.6,"Región de Murcia"
"Y15-24","ES63",2007,38.3,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2007,31.5,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2007,22.1,"Canarias (ES)"
"Y15-24","ES70",2007,22.1,"Canarias (ES)"
"Y15-24","EU15",2007,15,"European Union (15 countries)"
"Y15-24","EU27",2007,15.6,"European Union (27 countries)"
"Y15-24","EU28",2007,15.6,"European Union (28 countries)"
"Y15-24","FI",2007,16.5,"Finland"
"Y15-24","FI1",2007,16.5,"Manner-Suomi"
"Y15-24","FI19",2007,14.9,"Länsi-Suomi"
"Y15-24","FI1B",2007,13,"Helsinki-Uusimaa"
"Y15-24","FI1C",2007,16.4,"Etelä-Suomi"
"Y15-24","FI1D",2007,22.9,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2007,NA,"Åland"
"Y15-24","FI20",2007,NA,"Åland"
"Y15-24","FR",2007,19.5,"France"
"Y15-24","FR1",2007,17.8,"Île de France"
"Y15-24","FR10",2007,17.8,"Île de France"
"Y15-24","FR2",2007,19.3,"Bassin Parisien"
"Y15-24","FR21",2007,20.7,"Champagne-Ardenne"
"Y15-24","FR22",2007,22.9,"Picardie"
"Y15-24","FR23",2007,22.8,"Haute-Normandie"
"Y15-24","FR24",2007,15.5,"Centre (FR)"
"Y15-24","FR25",2007,15,"Basse-Normandie"
"Y15-24","FR26",2007,15.9,"Bourgogne"
"Y15-24","FR3",2007,28.3,"Nord - Pas-de-Calais"
"Y15-24","FR30",2007,28.3,"Nord - Pas-de-Calais"
"Y15-24","FR4",2007,16.8,"Est (FR)"
"Y15-24","FR41",2007,16.5,"Lorraine"
"Y15-24","FR42",2007,16.4,"Alsace"
"Y15-24","FR43",2007,18.2,"Franche-Comté"
"Y15-24","FR5",2007,14.3,"Ouest (FR)"
"Y15-24","FR51",2007,12.3,"Pays de la Loire"
"Y15-24","FR52",2007,14.1,"Bretagne"
"Y15-24","FR53",2007,19.4,"Poitou-Charentes"
"Y15-24","FR6",2007,20.2,"Sud-Ouest (FR)"
"Y15-24","FR61",2007,20.1,"Aquitaine"
"Y15-24","FR62",2007,21.3,"Midi-Pyrénées"
"Y15-24","FR63",2007,NA,"Limousin"
"Y15-24","FR7",2007,16.5,"Centre-Est (FR)"
"Y15-24","FR71",2007,15.9,"Rhône-Alpes"
"Y15-24","FR72",2007,19.3,"Auvergne"
"Y15-24","FR8",2007,22,"Méditerranée"
"Y15-24","FR81",2007,26,"Languedoc-Roussillon"
"Y15-24","FR82",2007,19.6,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2007,NA,"Corse"
"Y15-24","FR9",2007,46.9,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2007,53.3,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2007,45,"Martinique (NUTS 2010)"
"Y15-24","FR93",2007,39.9,"Guyane (NUTS 2010)"
"Y15-24","FR94",2007,46.8,"Réunion (NUTS 2010)"
"Y15-24","HR",2007,25.2,"Croatia"
"Y15-24","HR0",2007,25.2,"Hrvatska"
"Y15-24","HR03",2007,21.5,"Jadranska Hrvatska"
"Y15-24","HR04",2007,26.7,"Kontinentalna Hrvatska"
"Y15-24","HU",2007,18,"Hungary"
"Y15-24","HU1",2007,10.3,"Közép-Magyarország"
"Y15-24","HU10",2007,10.3,"Közép-Magyarország"
"Y15-24","HU2",2007,14.8,"Dunántúl"
"Y15-24","HU21",2007,11.4,"Közép-Dunántúl"
"Y15-24","HU22",2007,12,"Nyugat-Dunántúl"
"Y15-24","HU23",2007,23.4,"Dél-Dunántúl"
"Y15-24","HU3",2007,24.9,"Alföld és Észak"
"Y15-24","HU31",2007,27.6,"Észak-Magyarország"
"Y15-24","HU32",2007,26.8,"Észak-Alföld"
"Y15-24","HU33",2007,19.8,"Dél-Alföld"
"Y15-24","IE",2007,9.1,"Ireland"
"Y15-24","IE0",2007,9.1,"Éire/Ireland"
"Y15-24","IE01",2007,9.7,"Border, Midland and Western"
"Y15-24","IE02",2007,8.8,"Southern and Eastern"
"Y15-24","IS",2007,7,"Iceland"
"Y15-24","IS0",2007,7,"Ísland"
"Y15-24","IS00",2007,7,"Ísland"
"Y15-24","IT",2007,20.4,"Italy"
"Y15-24","ITC",2007,13.8,"Nord-Ovest"
"Y15-24","ITC1",2007,14.5,"Piemonte"
"Y15-24","ITC2",2007,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2007,19.9,"Liguria"
"Y15-24","ITC4",2007,12.9,"Lombardia"
"Y15-24","ITF",2007,30.5,"Sud"
"Y15-24","ITF1",2007,17.1,"Abruzzo"
"Y15-24","ITF2",2007,23.2,"Molise"
"Y15-24","ITF3",2007,32.5,"Campania"
"Y15-24","ITF4",2007,31.7,"Puglia"
"Y15-24","ITF5",2007,30.8,"Basilicata"
"Y15-24","ITF6",2007,31.2,"Calabria"
"Y15-24","ITG",2007,36.2,"Isole"
"Y15-24","ITG1",2007,37.7,"Sicilia"
"Y15-24","ITG2",2007,32,"Sardegna"
"Y15-24","ITH",2007,9.6,"Nord-Est"
"Y15-24","ITH1",2007,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2007,9.1,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2007,8.5,"Veneto"
"Y15-24","ITH4",2007,14.5,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2007,10.7,"Emilia-Romagna"
"Y15-24","ITI",2007,18,"Centro (IT)"
"Y15-24","ITI1",2007,13.9,"Toscana"
"Y15-24","ITI2",2007,12.8,"Umbria"
"Y15-24","ITI3",2007,8.9,"Marche"
"Y15-24","ITI4",2007,25.6,"Lazio"
"Y15-24","LT",2007,8.4,"Lithuania"
"Y15-24","LT0",2007,8.4,"Lietuva"
"Y15-24","LT00",2007,8.4,"Lietuva"
"Y15-24","LU",2007,15.2,"Luxembourg"
"Y15-24","LU0",2007,15.2,"Luxembourg"
"Y15-24","LU00",2007,15.2,"Luxembourg"
"Y15-24","LV",2007,10.6,"Latvia"
"Y15-24","LV0",2007,10.6,"Latvija"
"Y15-24","LV00",2007,10.6,"Latvija"
"Y15-24","MK",2007,57.7,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2007,57.7,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2007,57.7,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2007,13.5,"Malta"
"Y15-24","MT0",2007,13.5,"Malta"
"Y15-24","MT00",2007,13.5,"Malta"
"Y15-24","NL",2007,5.9,"Netherlands"
"Y15-24","NL1",2007,7.6,"Noord-Nederland"
"Y15-24","NL11",2007,8.9,"Groningen"
"Y15-24","NL12",2007,6,"Friesland (NL)"
"Y15-24","NL13",2007,7.9,"Drenthe"
"Y15-24","NL2",2007,5.2,"Oost-Nederland"
"Y15-24","NL21",2007,5.1,"Overijssel"
"Y15-24","NL22",2007,4.9,"Gelderland"
"Y15-24","NL23",2007,7,"Flevoland"
"Y15-24","NL3",2007,5.9,"West-Nederland"
"Y15-24","NL31",2007,5,"Utrecht"
"Y15-24","NL32",2007,5.6,"Noord-Holland"
"Y15-24","NL33",2007,6.6,"Zuid-Holland"
"Y15-24","NL34",2007,5.2,"Zeeland"
"Y15-24","NL4",2007,5.9,"Zuid-Nederland"
"Y15-24","NL41",2007,5.2,"Noord-Brabant"
"Y15-24","NL42",2007,7.4,"Limburg (NL)"
"Y15-24","NO",2007,7.4,"Norway"
"Y15-24","NO0",2007,7.4,"Norge"
"Y15-24","NO01",2007,7.8,"Oslo og Akershus"
"Y15-24","NO02",2007,9.1,"Hedmark og Oppland"
"Y15-24","NO03",2007,7.7,"Sør-Østlandet"
"Y15-24","NO04",2007,5.1,"Agder og Rogaland"
"Y15-24","NO05",2007,6.7,"Vestlandet"
"Y15-24","NO06",2007,9.4,"Trøndelag"
"Y15-24","NO07",2007,8.3,"Nord-Norge"
"Y15-24","PL",2007,21.7,"Poland"
"Y15-24","PL1",2007,20.1,"Region Centralny"
"Y15-24","PL11",2007,17.8,"Lódzkie"
"Y15-24","PL12",2007,21.3,"Mazowieckie"
"Y15-24","PL2",2007,20.6,"Region Poludniowy"
"Y15-24","PL21",2007,24.2,"Malopolskie"
"Y15-24","PL22",2007,17.5,"Slaskie"
"Y15-24","PL3",2007,24.3,"Region Wschodni"
"Y15-24","PL31",2007,24.3,"Lubelskie"
"Y15-24","PL32",2007,24.4,"Podkarpackie"
"Y15-24","PL33",2007,27.8,"Swietokrzyskie"
"Y15-24","PL34",2007,19.7,"Podlaskie"
"Y15-24","PL4",2007,21.2,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2007,19.3,"Wielkopolskie"
"Y15-24","PL42",2007,24.5,"Zachodniopomorskie"
"Y15-24","PL43",2007,25.1,"Lubuskie"
"Y15-24","PL5",2007,21.7,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2007,22.8,"Dolnoslaskie"
"Y15-24","PL52",2007,18.3,"Opolskie"
"Y15-24","PL6",2007,22.6,"Region Pólnocny"
"Y15-24","PL61",2007,22.9,"Kujawsko-Pomorskie"
"Y15-24","PL62",2007,25.1,"Warminsko-Mazurskie"
"Y15-24","PL63",2007,20.8,"Pomorskie"
"Y15-24","PT",2007,16.7,"Portugal"
"Y15-24","PT1",2007,16.9,"Continente"
"Y15-24","PT11",2007,16.8,"Norte"
"Y15-24","PT15",2007,NA,"Algarve"
"Y15-24","PT16",2007,13.7,"Centro (PT)"
"Y15-24","PT17",2007,18.6,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2007,20.3,"Alentejo"
"Y15-24","PT2",2007,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2007,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2007,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2007,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2007,20.1,"Romania"
"Y15-24","RO1",2007,19.4,"Macroregiunea unu"
"Y15-24","RO11",2007,14.1,"Nord-Vest"
"Y15-24","RO12",2007,24.7,"Centru"
"Y15-24","RO2",2007,19.7,"Macroregiunea doi"
"Y15-24","RO21",2007,14.7,"Nord-Est"
"Y15-24","RO22",2007,26.5,"Sud-Est"
"Y15-24","RO3",2007,21.6,"Macroregiunea trei"
"Y15-24","RO31",2007,23.9,"Sud - Muntenia"
"Y15-24","RO32",2007,16.1,"Bucuresti - Ilfov"
"Y15-24","RO4",2007,19.8,"Macroregiunea patru"
"Y15-24","RO41",2007,22.1,"Sud-Vest Oltenia"
"Y15-24","RO42",2007,17.3,"Vest"
"Y15-24","SE",2007,19.3,"Sweden"
"Y15-24","SE1",2007,20.2,"Östra Sverige"
"Y15-24","SE11",2007,20.1,"Stockholm"
"Y15-24","SE12",2007,20.2,"Östra Mellansverige"
"Y15-24","SE2",2007,18.7,"Södra Sverige"
"Y15-24","SE21",2007,15.8,"Småland med öarna"
"Y15-24","SE22",2007,22.1,"Sydsverige"
"Y15-24","SE23",2007,17.7,"Västsverige"
"Y15-24","SE3",2007,19.1,"Norra Sverige"
"Y15-24","SE31",2007,18.7,"Norra Mellansverige"
"Y15-24","SE32",2007,20,"Mellersta Norrland"
"Y15-24","SE33",2007,19.2,"Övre Norrland"
"Y15-24","SI",2007,10.1,"Slovenia"
"Y15-24","SI0",2007,10.1,"Slovenija"
"Y15-24","SI01",2007,12.3,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2007,7.6,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2007,20.3,"Slovakia"
"Y15-24","SK0",2007,20.3,"Slovensko"
"Y15-24","SK01",2007,7.6,"Bratislavský kraj"
"Y15-24","SK02",2007,13,"Západné Slovensko"
"Y15-24","SK03",2007,24.7,"Stredné Slovensko"
"Y15-24","SK04",2007,29.6,"Východné Slovensko"
"Y15-24","TR",2007,17.2,"Turkey"
"Y15-24","TR1",2007,15.5,"Istanbul"
"Y15-24","TR10",2007,15.5,"Istanbul"
"Y15-24","TR2",2007,13.3,"Bati Marmara"
"Y15-24","TR21",2007,15.6,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2007,10.8,"Balikesir, Çanakkale"
"Y15-24","TR3",2007,14.3,"Ege"
"Y15-24","TR31",2007,17.1,"Izmir"
"Y15-24","TR32",2007,14.2,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2007,10.4,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2007,17.8,"Dogu Marmara"
"Y15-24","TR41",2007,15,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2007,21.4,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2007,22.2,"Bati Anadolu"
"Y15-24","TR51",2007,25.2,"Ankara"
"Y15-24","TR52",2007,17.1,"Konya, Karaman"
"Y15-24","TR6",2007,18.1,"Akdeniz"
"Y15-24","TR61",2007,11.5,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2007,23.6,"Adana, Mersin"
"Y15-24","TR63",2007,17.7,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2007,20.5,"Orta Anadolu"
"Y15-24","TR71",2007,17.3,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2007,22.6,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2007,14.5,"Bati Karadeniz"
"Y15-24","TR81",2007,19.3,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2007,7.7,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2007,14.4,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2007,15.5,"Dogu Karadeniz"
"Y15-24","TR90",2007,15.5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2007,7.9,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2007,8.4,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2007,7.5,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2007,22.9,"Ortadogu Anadolu"
"Y15-24","TRB1",2007,28,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2007,19.2,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2007,23,"Güneydogu Anadolu"
"Y15-24","TRC1",2007,22,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2007,21.2,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2007,28.4,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2007,14.3,"United Kingdom"
"Y15-24","UKC",2007,16,"North East (UK)"
"Y15-24","UKC1",2007,17.7,"Tees Valley and Durham"
"Y15-24","UKC2",2007,14.8,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2007,15.1,"North West (UK)"
"Y15-24","UKD1",2007,NA,"Cumbria"
"Y15-24","UKD3",2007,15.6,"Greater Manchester"
"Y15-24","UKD4",2007,13.6,"Lancashire"
"Y15-24","UKD6",2007,9.8,"Cheshire"
"Y15-24","UKD7",2007,20,"Merseyside"
"Y15-24","UKE",2007,14,"Yorkshire and The Humber"
"Y15-24","UKE1",2007,15.1,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2007,10.4,"North Yorkshire"
"Y15-24","UKE3",2007,14,"South Yorkshire"
"Y15-24","UKE4",2007,14.5,"West Yorkshire"
"Y15-24","UKF",2007,14.6,"East Midlands (UK)"
"Y15-24","UKF1",2007,16.4,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2007,13,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2007,13.9,"Lincolnshire"
"Y15-24","UKG",2007,16.9,"West Midlands (UK)"
"Y15-24","UKG1",2007,11.7,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2007,14.3,"Shropshire and Staffordshire"
"Y15-24","UKG3",2007,20.5,"West Midlands"
"Y15-24","UKH",2007,12.7,"East of England"
"Y15-24","UKH1",2007,12.1,"East Anglia"
"Y15-24","UKH2",2007,14.2,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2007,12.4,"Essex"
"Y15-24","UKI",2007,18.4,"London"
"Y15-24","UKI1",2007,21.2,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2007,16.7,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2007,12.7,"South East (UK)"
"Y15-24","UKJ1",2007,11.6,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2007,12.2,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2007,11.7,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2007,15.7,"Kent"
"Y15-24","UKK",2007,10.6,"South West (UK)"
"Y15-24","UKK1",2007,8.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2007,11,"Dorset and Somerset"
"Y15-24","UKK3",2007,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2007,13.8,"Devon"
"Y15-24","UKL",2007,14.5,"Wales"
"Y15-24","UKL1",2007,14.7,"West Wales and The Valleys"
"Y15-24","UKL2",2007,14.1,"East Wales"
"Y15-24","UKM",2007,13.2,"Scotland"
"Y15-24","UKM2",2007,15.4,"Eastern Scotland"
"Y15-24","UKM3",2007,13.4,"South Western Scotland"
"Y15-24","UKM5",2007,NA,"North Eastern Scotland"
"Y15-24","UKM6",2007,NA,"Highlands and Islands"
"Y15-24","UKN",2007,9.3,"Northern Ireland (UK)"
"Y15-24","UKN0",2007,9.3,"Northern Ireland (UK)"
"Y20-64","AT",2007,4.5,"Austria"
"Y20-64","AT1",2007,6.1,"Ostösterreich"
"Y20-64","AT11",2007,3.8,"Burgenland (AT)"
"Y20-64","AT12",2007,3.7,"Niederösterreich"
"Y20-64","AT13",2007,8.7,"Wien"
"Y20-64","AT2",2007,3.8,"Südösterreich"
"Y20-64","AT21",2007,3.9,"Kärnten"
"Y20-64","AT22",2007,3.7,"Steiermark"
"Y20-64","AT3",2007,3.2,"Westösterreich"
"Y20-64","AT31",2007,3.2,"Oberösterreich"
"Y20-64","AT32",2007,3.3,"Salzburg"
"Y20-64","AT33",2007,2.7,"Tirol"
"Y20-64","AT34",2007,3.7,"Vorarlberg"
"Y20-64","BE",2007,7.2,"Belgium"
"Y20-64","BE1",2007,16.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2007,16.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2007,4.1,"Vlaams Gewest"
"Y20-64","BE21",2007,4.7,"Prov. Antwerpen"
"Y20-64","BE22",2007,5.1,"Prov. Limburg (BE)"
"Y20-64","BE23",2007,4.6,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2007,3.2,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2007,2.8,"Prov. West-Vlaanderen"
"Y20-64","BE3",2007,10.2,"Région wallonne"
"Y20-64","BE31",2007,6.9,"Prov. Brabant Wallon"
"Y20-64","BE32",2007,12.3,"Prov. Hainaut"
"Y20-64","BE33",2007,10.6,"Prov. Liège"
"Y20-64","BE34",2007,6.4,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2007,8.2,"Prov. Namur"
"Y20-64","BG",2007,6.6,"Bulgaria"
"Y20-64","BG3",2007,8.9,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2007,8.6,"Severozapaden"
"Y20-64","BG32",2007,10.2,"Severen tsentralen"
"Y20-64","BG33",2007,10.5,"Severoiztochen"
"Y20-64","BG34",2007,6.3,"Yugoiztochen"
"Y20-64","BG4",2007,4.5,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2007,3.8,"Yugozapaden"
"Y20-64","BG42",2007,5.5,"Yuzhen tsentralen"
"Y20-64","CH",2007,3.5,"Switzerland"
"Y20-64","CH0",2007,3.5,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2007,4.5,"Région lémanique"
"Y20-64","CH02",2007,4,"Espace Mittelland"
"Y20-64","CH03",2007,3,"Nordwestschweiz"
"Y20-64","CH04",2007,3.4,"Zürich"
"Y20-64","CH05",2007,2.3,"Ostschweiz"
"Y20-64","CH06",2007,2.7,"Zentralschweiz"
"Y20-64","CH07",2007,5.1,"Ticino"
"Y20-64","CY",2007,3.9,"Cyprus"
"Y20-64","CY0",2007,3.9,"Kypros"
"Y20-64","CY00",2007,3.9,"Kypros"
"Y20-64","CZ",2007,5.2,"Czech Republic"
"Y20-64","CZ0",2007,5.2,"Ceská republika"
"Y20-64","CZ01",2007,2.4,"Praha"
"Y20-64","CZ02",2007,3.3,"Strední Cechy"
"Y20-64","CZ03",2007,3.3,"Jihozápad"
"Y20-64","CZ04",2007,9.1,"Severozápad"
"Y20-64","CZ05",2007,4.6,"Severovýchod"
"Y20-64","CZ06",2007,5.1,"Jihovýchod"
"Y20-64","CZ07",2007,5.9,"Strední Morava"
"Y20-64","CZ08",2007,8.3,"Moravskoslezsko"
"Y20-64","DE",2007,8.6,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2007,4.9,"Baden-Württemberg"
"Y20-64","DE11",2007,5,"Stuttgart"
"Y20-64","DE12",2007,5.4,"Karlsruhe"
"Y20-64","DE13",2007,4.3,"Freiburg"
"Y20-64","DE14",2007,4.6,"Tübingen"
"Y20-64","DE2",2007,5.2,"Bayern"
"Y20-64","DE21",2007,4.3,"Oberbayern"
"Y20-64","DE22",2007,5,"Niederbayern"
"Y20-64","DE23",2007,5.2,"Oberpfalz"
"Y20-64","DE24",2007,7.3,"Oberfranken"
"Y20-64","DE25",2007,6.5,"Mittelfranken"
"Y20-64","DE26",2007,5.4,"Unterfranken"
"Y20-64","DE27",2007,4.9,"Schwaben"
"Y20-64","DE3",2007,16.4,"Berlin"
"Y20-64","DE30",2007,16.4,"Berlin"
"Y20-64","DE4",2007,13.8,"Brandenburg"
"Y20-64","DE40",2007,13.8,"Brandenburg"
"Y20-64","DE5",2007,11.8,"Bremen"
"Y20-64","DE50",2007,11.8,"Bremen"
"Y20-64","DE6",2007,8.8,"Hamburg"
"Y20-64","DE60",2007,8.8,"Hamburg"
"Y20-64","DE7",2007,7.2,"Hessen"
"Y20-64","DE71",2007,7.1,"Darmstadt"
"Y20-64","DE72",2007,7,"Gießen"
"Y20-64","DE73",2007,7.8,"Kassel"
"Y20-64","DE8",2007,17.8,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2007,17.8,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2007,7.8,"Niedersachsen"
"Y20-64","DE91",2007,8.8,"Braunschweig"
"Y20-64","DE92",2007,8.5,"Hannover"
"Y20-64","DE93",2007,7.4,"Lüneburg"
"Y20-64","DE94",2007,7,"Weser-Ems"
"Y20-64","DEA",2007,8.2,"Nordrhein-Westfalen"
"Y20-64","DEA1",2007,8.4,"Düsseldorf"
"Y20-64","DEA2",2007,7.7,"Köln"
"Y20-64","DEA3",2007,7.2,"Münster"
"Y20-64","DEA4",2007,8,"Detmold"
"Y20-64","DEA5",2007,9.5,"Arnsberg"
"Y20-64","DEB",2007,5.8,"Rheinland-Pfalz"
"Y20-64","DEB1",2007,6.1,"Koblenz"
"Y20-64","DEB2",2007,5.2,"Trier"
"Y20-64","DEB3",2007,5.7,"Rheinhessen-Pfalz"
"Y20-64","DEC",2007,7.1,"Saarland"
"Y20-64","DEC0",2007,7.1,"Saarland"
"Y20-64","DED",2007,14.7,"Sachsen"
"Y20-64","DED2",2007,13.5,"Dresden"
"Y20-64","DED4",2007,14.2,"Chemnitz"
"Y20-64","DED5",2007,17.4,"Leipzig"
"Y20-64","DEE",2007,15.6,"Sachsen-Anhalt"
"Y20-64","DEE0",2007,15.6,"Sachsen-Anhalt"
"Y20-64","DEF",2007,7.7,"Schleswig-Holstein"
"Y20-64","DEF0",2007,7.7,"Schleswig-Holstein"
"Y20-64","DEG",2007,13.9,"Thüringen"
"Y20-64","DEG0",2007,13.9,"Thüringen"
"Y20-64","DK",2007,3.4,"Denmark"
"Y20-64","DK0",2007,3.4,"Danmark"
"Y20-64","DK01",2007,4,"Hovedstaden"
"Y20-64","DK02",2007,3.2,"Sjælland"
"Y20-64","DK03",2007,3,"Syddanmark"
"Y20-64","DK04",2007,3,"Midtjylland"
"Y20-64","DK05",2007,4,"Nordjylland"
"Y20-64","EA17",2007,7.2,"Euro area (17 countries)"
"Y20-64","EA18",2007,7.2,"Euro area (18 countries)"
"Y20-64","EA19",2007,7.2,"Euro area (19 countries)"
"Y20-64","EE",2007,4.4,"Estonia"
"Y20-64","EE0",2007,4.4,"Eesti"
"Y20-64","EE00",2007,4.4,"Eesti"
"Y20-64","EL",2007,8.3,"Greece"
"Y20-64","EL1",2007,9.1,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2007,9.6,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2007,9,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2007,12.2,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2007,7.9,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2007,9,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2007,10,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2007,8.9,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2007,9.7,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2007,9.3,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2007,7.5,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2007,7.7,"Attiki"
"Y20-64","EL30",2007,7.7,"Attiki"
"Y20-64","EL4",2007,6.9,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2007,7.8,"Voreio Aigaio"
"Y20-64","EL42",2007,9.3,"Notio Aigaio"
"Y20-64","EL43",2007,5.5,"Kriti"
"Y20-64","ES",2007,7.8,"Spain"
"Y20-64","ES1",2007,7.3,"Noroeste (ES)"
"Y20-64","ES11",2007,7.3,"Galicia"
"Y20-64","ES12",2007,8.3,"Principado de Asturias"
"Y20-64","ES13",2007,5.8,"Cantabria"
"Y20-64","ES2",2007,5.4,"Noreste (ES)"
"Y20-64","ES21",2007,6,"País Vasco"
"Y20-64","ES22",2007,4.5,"Comunidad Foral de Navarra"
"Y20-64","ES23",2007,5.3,"La Rioja"
"Y20-64","ES24",2007,4.9,"Aragón"
"Y20-64","ES3",2007,5.8,"Comunidad de Madrid"
"Y20-64","ES30",2007,5.8,"Comunidad de Madrid"
"Y20-64","ES4",2007,7.9,"Centro (ES)"
"Y20-64","ES41",2007,6.8,"Castilla y León"
"Y20-64","ES42",2007,7.1,"Castilla-la Mancha"
"Y20-64","ES43",2007,12.5,"Extremadura"
"Y20-64","ES5",2007,6.9,"Este (ES)"
"Y20-64","ES51",2007,6.1,"Cataluña"
"Y20-64","ES52",2007,8.1,"Comunidad Valenciana"
"Y20-64","ES53",2007,6.8,"Illes Balears"
"Y20-64","ES6",2007,11.4,"Sur (ES)"
"Y20-64","ES61",2007,12.1,"Andalucía"
"Y20-64","ES62",2007,6.8,"Región de Murcia"
"Y20-64","ES63",2007,19.8,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2007,17.3,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2007,9.9,"Canarias (ES)"
"Y20-64","ES70",2007,9.9,"Canarias (ES)"
"Y20-64","EU15",2007,6.7,"European Union (15 countries)"
"Y20-64","EU27",2007,6.8,"European Union (27 countries)"
"Y20-64","EU28",2007,6.9,"European Union (28 countries)"
"Y20-64","FI",2007,6.1,"Finland"
"Y20-64","FI1",2007,6.2,"Manner-Suomi"
"Y20-64","FI19",2007,5.9,"Länsi-Suomi"
"Y20-64","FI1B",2007,4.3,"Helsinki-Uusimaa"
"Y20-64","FI1C",2007,6,"Etelä-Suomi"
"Y20-64","FI1D",2007,9.1,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2007,NA,"Åland"
"Y20-64","FI20",2007,NA,"Åland"
"Y20-64","FR",2007,7.6,"France"
"Y20-64","FR1",2007,7.5,"Île de France"
"Y20-64","FR10",2007,7.5,"Île de France"
"Y20-64","FR2",2007,6.9,"Bassin Parisien"
"Y20-64","FR21",2007,7.5,"Champagne-Ardenne"
"Y20-64","FR22",2007,9.3,"Picardie"
"Y20-64","FR23",2007,7.8,"Haute-Normandie"
"Y20-64","FR24",2007,5.3,"Centre (FR)"
"Y20-64","FR25",2007,5.3,"Basse-Normandie"
"Y20-64","FR26",2007,6.5,"Bourgogne"
"Y20-64","FR3",2007,10.7,"Nord - Pas-de-Calais"
"Y20-64","FR30",2007,10.7,"Nord - Pas-de-Calais"
"Y20-64","FR4",2007,6.5,"Est (FR)"
"Y20-64","FR41",2007,7,"Lorraine"
"Y20-64","FR42",2007,5.6,"Alsace"
"Y20-64","FR43",2007,6.8,"Franche-Comté"
"Y20-64","FR5",2007,6,"Ouest (FR)"
"Y20-64","FR51",2007,5.6,"Pays de la Loire"
"Y20-64","FR52",2007,6.5,"Bretagne"
"Y20-64","FR53",2007,5.8,"Poitou-Charentes"
"Y20-64","FR6",2007,6.9,"Sud-Ouest (FR)"
"Y20-64","FR61",2007,6.4,"Aquitaine"
"Y20-64","FR62",2007,7.5,"Midi-Pyrénées"
"Y20-64","FR63",2007,6.3,"Limousin"
"Y20-64","FR7",2007,6.3,"Centre-Est (FR)"
"Y20-64","FR71",2007,6,"Rhône-Alpes"
"Y20-64","FR72",2007,7.8,"Auvergne"
"Y20-64","FR8",2007,9,"Méditerranée"
"Y20-64","FR81",2007,9.7,"Languedoc-Roussillon"
"Y20-64","FR82",2007,8.6,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2007,11.4,"Corse"
"Y20-64","FR9",2007,21.8,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2007,22.4,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2007,20.5,"Martinique (NUTS 2010)"
"Y20-64","FR93",2007,19.8,"Guyane (NUTS 2010)"
"Y20-64","FR94",2007,22.7,"Réunion (NUTS 2010)"
"Y20-64","HR",2007,9.4,"Croatia"
"Y20-64","HR0",2007,9.4,"Hrvatska"
"Y20-64","HR03",2007,8.7,"Jadranska Hrvatska"
"Y20-64","HR04",2007,9.8,"Kontinentalna Hrvatska"
"Y20-64","HU",2007,7.3,"Hungary"
"Y20-64","HU1",2007,4.7,"Közép-Magyarország"
"Y20-64","HU10",2007,4.7,"Közép-Magyarország"
"Y20-64","HU2",2007,6.3,"Dunántúl"
"Y20-64","HU21",2007,4.8,"Közép-Dunántúl"
"Y20-64","HU22",2007,5,"Nyugat-Dunántúl"
"Y20-64","HU23",2007,9.8,"Dél-Dunántúl"
"Y20-64","HU3",2007,10.1,"Alföld és Észak"
"Y20-64","HU31",2007,12.3,"Észak-Magyarország"
"Y20-64","HU32",2007,10.5,"Észak-Alföld"
"Y20-64","HU33",2007,7.9,"Dél-Alföld"
"Y20-64","IE",2007,4.4,"Ireland"
"Y20-64","IE0",2007,4.4,"Éire/Ireland"
"Y20-64","IE01",2007,4.7,"Border, Midland and Western"
"Y20-64","IE02",2007,4.3,"Southern and Eastern"
"Y20-64","IS",2007,1.6,"Iceland"
"Y20-64","IS0",2007,1.6,"Ísland"
"Y20-64","IS00",2007,1.6,"Ísland"
"Y20-64","IT",2007,5.8,"Italy"
"Y20-64","ITC",2007,3.5,"Nord-Ovest"
"Y20-64","ITC1",2007,4,"Piemonte"
"Y20-64","ITC2",2007,2.9,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2007,4.6,"Liguria"
"Y20-64","ITC4",2007,3.1,"Lombardia"
"Y20-64","ITF",2007,10,"Sud"
"Y20-64","ITF1",2007,6.1,"Abruzzo"
"Y20-64","ITF2",2007,7.8,"Molise"
"Y20-64","ITF3",2007,10.8,"Campania"
"Y20-64","ITF4",2007,10.5,"Puglia"
"Y20-64","ITF5",2007,9.2,"Basilicata"
"Y20-64","ITF6",2007,10.8,"Calabria"
"Y20-64","ITG",2007,11.5,"Isole"
"Y20-64","ITG1",2007,12.3,"Sicilia"
"Y20-64","ITG2",2007,9.5,"Sardegna"
"Y20-64","ITH",2007,3,"Nord-Est"
"Y20-64","ITH1",2007,2.5,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2007,2.7,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2007,3.2,"Veneto"
"Y20-64","ITH4",2007,3.2,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2007,2.7,"Emilia-Romagna"
"Y20-64","ITI",2007,5.1,"Centro (IT)"
"Y20-64","ITI1",2007,4.2,"Toscana"
"Y20-64","ITI2",2007,4.6,"Umbria"
"Y20-64","ITI3",2007,4.1,"Marche"
"Y20-64","ITI4",2007,6.2,"Lazio"
"Y20-64","LT",2007,4.2,"Lithuania"
"Y20-64","LT0",2007,4.2,"Lietuva"
"Y20-64","LT00",2007,4.2,"Lietuva"
"Y20-64","LU",2007,3.8,"Luxembourg"
"Y20-64","LU0",2007,3.8,"Luxembourg"
"Y20-64","LU00",2007,3.8,"Luxembourg"
"Y20-64","LV",2007,5.8,"Latvia"
"Y20-64","LV0",2007,5.8,"Latvija"
"Y20-64","LV00",2007,5.8,"Latvija"
"Y20-64","MK",2007,34.3,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2007,34.3,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2007,34.3,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2007,5.4,"Malta"
"Y20-64","MT0",2007,5.4,"Malta"
"Y20-64","MT00",2007,5.4,"Malta"
"Y20-64","NL",2007,2.8,"Netherlands"
"Y20-64","NL1",2007,3.5,"Noord-Nederland"
"Y20-64","NL11",2007,4.4,"Groningen"
"Y20-64","NL12",2007,2.7,"Friesland (NL)"
"Y20-64","NL13",2007,3.3,"Drenthe"
"Y20-64","NL2",2007,2.7,"Oost-Nederland"
"Y20-64","NL21",2007,2.9,"Overijssel"
"Y20-64","NL22",2007,2.4,"Gelderland"
"Y20-64","NL23",2007,3.6,"Flevoland"
"Y20-64","NL3",2007,2.7,"West-Nederland"
"Y20-64","NL31",2007,2.2,"Utrecht"
"Y20-64","NL32",2007,2.6,"Noord-Holland"
"Y20-64","NL33",2007,3,"Zuid-Holland"
"Y20-64","NL34",2007,1.8,"Zeeland"
"Y20-64","NL4",2007,2.7,"Zuid-Nederland"
"Y20-64","NL41",2007,2.4,"Noord-Brabant"
"Y20-64","NL42",2007,3.5,"Limburg (NL)"
"Y20-64","NO",2007,2.1,"Norway"
"Y20-64","NO0",2007,2.1,"Norge"
"Y20-64","NO01",2007,2,"Oslo og Akershus"
"Y20-64","NO02",2007,1.8,"Hedmark og Oppland"
"Y20-64","NO03",2007,2.4,"Sør-Østlandet"
"Y20-64","NO04",2007,1.6,"Agder og Rogaland"
"Y20-64","NO05",2007,1.8,"Vestlandet"
"Y20-64","NO06",2007,2.6,"Trøndelag"
"Y20-64","NO07",2007,2.1,"Nord-Norge"
"Y20-64","PL",2007,9.6,"Poland"
"Y20-64","PL1",2007,9.1,"Region Centralny"
"Y20-64","PL11",2007,9.3,"Lódzkie"
"Y20-64","PL12",2007,8.9,"Mazowieckie"
"Y20-64","PL2",2007,8.1,"Region Poludniowy"
"Y20-64","PL21",2007,8.3,"Malopolskie"
"Y20-64","PL22",2007,8,"Slaskie"
"Y20-64","PL3",2007,10.1,"Region Wschodni"
"Y20-64","PL31",2007,9.7,"Lubelskie"
"Y20-64","PL32",2007,9.7,"Podkarpackie"
"Y20-64","PL33",2007,12.1,"Swietokrzyskie"
"Y20-64","PL34",2007,9,"Podlaskie"
"Y20-64","PL4",2007,9.3,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2007,8.2,"Wielkopolskie"
"Y20-64","PL42",2007,11.4,"Zachodniopomorskie"
"Y20-64","PL43",2007,9.7,"Lubuskie"
"Y20-64","PL5",2007,11.8,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2007,12.6,"Dolnoslaskie"
"Y20-64","PL52",2007,9.4,"Opolskie"
"Y20-64","PL6",2007,10.3,"Region Pólnocny"
"Y20-64","PL61",2007,11.3,"Kujawsko-Pomorskie"
"Y20-64","PL62",2007,10.2,"Warminsko-Mazurskie"
"Y20-64","PL63",2007,9.4,"Pomorskie"
"Y20-64","PT",2007,8.2,"Portugal"
"Y20-64","PT1",2007,8.3,"Continente"
"Y20-64","PT11",2007,9.5,"Norte"
"Y20-64","PT15",2007,6.5,"Algarve"
"Y20-64","PT16",2007,6.2,"Centro (PT)"
"Y20-64","PT17",2007,8.8,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2007,8.3,"Alentejo"
"Y20-64","PT2",2007,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2007,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2007,6.6,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2007,6.6,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2007,6.3,"Romania"
"Y20-64","RO1",2007,6,"Macroregiunea unu"
"Y20-64","RO11",2007,4,"Nord-Vest"
"Y20-64","RO12",2007,8.1,"Centru"
"Y20-64","RO2",2007,6.4,"Macroregiunea doi"
"Y20-64","RO21",2007,5,"Nord-Est"
"Y20-64","RO22",2007,8.2,"Sud-Est"
"Y20-64","RO3",2007,6.4,"Macroregiunea trei"
"Y20-64","RO31",2007,8.2,"Sud - Muntenia"
"Y20-64","RO32",2007,3.8,"Bucuresti - Ilfov"
"Y20-64","RO4",2007,6.3,"Macroregiunea patru"
"Y20-64","RO41",2007,7.2,"Sud-Vest Oltenia"
"Y20-64","RO42",2007,5.2,"Vest"
"Y20-64","SE",2007,5.1,"Sweden"
"Y20-64","SE1",2007,5.1,"Östra Sverige"
"Y20-64","SE11",2007,4.6,"Stockholm"
"Y20-64","SE12",2007,5.8,"Östra Mellansverige"
"Y20-64","SE2",2007,5,"Södra Sverige"
"Y20-64","SE21",2007,4.3,"Småland med öarna"
"Y20-64","SE22",2007,5.7,"Sydsverige"
"Y20-64","SE23",2007,4.8,"Västsverige"
"Y20-64","SE3",2007,5.5,"Norra Sverige"
"Y20-64","SE31",2007,5.4,"Norra Mellansverige"
"Y20-64","SE32",2007,5.1,"Mellersta Norrland"
"Y20-64","SE33",2007,6,"Övre Norrland"
"Y20-64","SI",2007,4.8,"Slovenia"
"Y20-64","SI0",2007,4.8,"Slovenija"
"Y20-64","SI01",2007,5.7,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2007,3.9,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2007,10.7,"Slovakia"
"Y20-64","SK0",2007,10.7,"Slovensko"
"Y20-64","SK01",2007,4.2,"Bratislavský kraj"
"Y20-64","SK02",2007,7.6,"Západné Slovensko"
"Y20-64","SK03",2007,14.7,"Stredné Slovensko"
"Y20-64","SK04",2007,14.2,"Východné Slovensko"
"Y20-64","TR",2007,8.5,"Turkey"
"Y20-64","TR1",2007,8.8,"Istanbul"
"Y20-64","TR10",2007,8.8,"Istanbul"
"Y20-64","TR2",2007,5.4,"Bati Marmara"
"Y20-64","TR21",2007,6.2,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2007,4.6,"Balikesir, Çanakkale"
"Y20-64","TR3",2007,7.6,"Ege"
"Y20-64","TR31",2007,8.9,"Izmir"
"Y20-64","TR32",2007,7.9,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2007,5.4,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2007,8,"Dogu Marmara"
"Y20-64","TR41",2007,6.9,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2007,9.4,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2007,9.4,"Bati Anadolu"
"Y20-64","TR51",2007,9.8,"Ankara"
"Y20-64","TR52",2007,8.6,"Konya, Karaman"
"Y20-64","TR6",2007,9.6,"Akdeniz"
"Y20-64","TR61",2007,5.8,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2007,12.7,"Adana, Mersin"
"Y20-64","TR63",2007,9.6,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2007,8.2,"Orta Anadolu"
"Y20-64","TR71",2007,6.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2007,9,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2007,6.5,"Bati Karadeniz"
"Y20-64","TR81",2007,6.9,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2007,3.3,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2007,7.2,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2007,4.8,"Dogu Karadeniz"
"Y20-64","TR90",2007,4.8,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2007,4.3,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2007,4.2,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2007,4.3,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2007,10.4,"Ortadogu Anadolu"
"Y20-64","TRB1",2007,10.1,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2007,10.7,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2007,15,"Güneydogu Anadolu"
"Y20-64","TRC1",2007,16.5,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2007,11.6,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2007,17.7,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2007,4.4,"United Kingdom"
"Y20-64","UKC",2007,5,"North East (UK)"
"Y20-64","UKC1",2007,4.7,"Tees Valley and Durham"
"Y20-64","UKC2",2007,5.2,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2007,4.9,"North West (UK)"
"Y20-64","UKD1",2007,3.3,"Cumbria"
"Y20-64","UKD3",2007,5.3,"Greater Manchester"
"Y20-64","UKD4",2007,4.8,"Lancashire"
"Y20-64","UKD6",2007,2.3,"Cheshire"
"Y20-64","UKD7",2007,6.5,"Merseyside"
"Y20-64","UKE",2007,4.4,"Yorkshire and The Humber"
"Y20-64","UKE1",2007,4.9,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2007,2.7,"North Yorkshire"
"Y20-64","UKE3",2007,5,"South Yorkshire"
"Y20-64","UKE4",2007,4.4,"West Yorkshire"
"Y20-64","UKF",2007,4.2,"East Midlands (UK)"
"Y20-64","UKF1",2007,4.8,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2007,3.6,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2007,4,"Lincolnshire"
"Y20-64","UKG",2007,5.2,"West Midlands (UK)"
"Y20-64","UKG1",2007,3,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2007,4.2,"Shropshire and Staffordshire"
"Y20-64","UKG3",2007,6.9,"West Midlands"
"Y20-64","UKH",2007,3.9,"East of England"
"Y20-64","UKH1",2007,3.5,"East Anglia"
"Y20-64","UKH2",2007,3.9,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2007,4.4,"Essex"
"Y20-64","UKI",2007,6,"London"
"Y20-64","UKI1",2007,7.4,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2007,5,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2007,3.6,"South East (UK)"
"Y20-64","UKJ1",2007,3.4,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2007,3.2,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2007,3.5,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2007,4.4,"Kent"
"Y20-64","UKK",2007,3.2,"South West (UK)"
"Y20-64","UKK1",2007,2.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2007,3.1,"Dorset and Somerset"
"Y20-64","UKK3",2007,4,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2007,3.7,"Devon"
"Y20-64","UKL",2007,4.3,"Wales"
"Y20-64","UKL1",2007,4.6,"West Wales and The Valleys"
"Y20-64","UKL2",2007,4,"East Wales"
"Y20-64","UKM",2007,3.9,"Scotland"
"Y20-64","UKM2",2007,4.3,"Eastern Scotland"
"Y20-64","UKM3",2007,4.2,"South Western Scotland"
"Y20-64","UKM5",2007,2.7,"North Eastern Scotland"
"Y20-64","UKM6",2007,1.9,"Highlands and Islands"
"Y20-64","UKN",2007,3.3,"Northern Ireland (UK)"
"Y20-64","UKN0",2007,3.3,"Northern Ireland (UK)"
"Y_GE15","AT",2007,4.9,"Austria"
"Y_GE15","AT1",2007,6.5,"Ostösterreich"
"Y_GE15","AT11",2007,4.1,"Burgenland (AT)"
"Y_GE15","AT12",2007,4,"Niederösterreich"
"Y_GE15","AT13",2007,9.2,"Wien"
"Y_GE15","AT2",2007,4.2,"Südösterreich"
"Y_GE15","AT21",2007,4.2,"Kärnten"
"Y_GE15","AT22",2007,4.1,"Steiermark"
"Y_GE15","AT3",2007,3.4,"Westösterreich"
"Y_GE15","AT31",2007,3.4,"Oberösterreich"
"Y_GE15","AT32",2007,3.5,"Salzburg"
"Y_GE15","AT33",2007,3,"Tirol"
"Y_GE15","AT34",2007,4.1,"Vorarlberg"
"Y_GE15","BE",2007,7.5,"Belgium"
"Y_GE15","BE1",2007,17.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2007,17.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2007,4.3,"Vlaams Gewest"
"Y_GE15","BE21",2007,5,"Prov. Antwerpen"
"Y_GE15","BE22",2007,5.3,"Prov. Limburg (BE)"
"Y_GE15","BE23",2007,4.8,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2007,3.4,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2007,3,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2007,10.5,"Région wallonne"
"Y_GE15","BE31",2007,7,"Prov. Brabant Wallon"
"Y_GE15","BE32",2007,12.8,"Prov. Hainaut"
"Y_GE15","BE33",2007,10.9,"Prov. Liège"
"Y_GE15","BE34",2007,6.8,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2007,8.5,"Prov. Namur"
"Y_GE15","BG",2007,6.9,"Bulgaria"
"Y_GE15","BG3",2007,9.2,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2007,9,"Severozapaden"
"Y_GE15","BG32",2007,10.7,"Severen tsentralen"
"Y_GE15","BG33",2007,10.8,"Severoiztochen"
"Y_GE15","BG34",2007,6.5,"Yugoiztochen"
"Y_GE15","BG4",2007,4.6,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2007,3.9,"Yugozapaden"
"Y_GE15","BG42",2007,5.6,"Yuzhen tsentralen"
"Y_GE15","CH",2007,3.7,"Switzerland"
"Y_GE15","CH0",2007,3.7,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2007,4.8,"Région lémanique"
"Y_GE15","CH02",2007,4.1,"Espace Mittelland"
"Y_GE15","CH03",2007,3.1,"Nordwestschweiz"
"Y_GE15","CH04",2007,3.4,"Zürich"
"Y_GE15","CH05",2007,2.6,"Ostschweiz"
"Y_GE15","CH06",2007,2.7,"Zentralschweiz"
"Y_GE15","CH07",2007,5,"Ticino"
"Y_GE15","CY",2007,3.9,"Cyprus"
"Y_GE15","CY0",2007,3.9,"Kypros"
"Y_GE15","CY00",2007,3.9,"Kypros"
"Y_GE15","CZ",2007,5.3,"Czech Republic"
"Y_GE15","CZ0",2007,5.3,"Ceská republika"
"Y_GE15","CZ01",2007,2.4,"Praha"
"Y_GE15","CZ02",2007,3.4,"Strední Cechy"
"Y_GE15","CZ03",2007,3.5,"Jihozápad"
"Y_GE15","CZ04",2007,9.5,"Severozápad"
"Y_GE15","CZ05",2007,4.8,"Severovýchod"
"Y_GE15","CZ06",2007,5.2,"Jihovýchod"
"Y_GE15","CZ07",2007,5.9,"Strední Morava"
"Y_GE15","CZ08",2007,8.5,"Moravskoslezsko"
"Y_GE15","DE",2007,8.7,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2007,5,"Baden-Württemberg"
"Y_GE15","DE11",2007,5.1,"Stuttgart"
"Y_GE15","DE12",2007,5.5,"Karlsruhe"
"Y_GE15","DE13",2007,4.3,"Freiburg"
"Y_GE15","DE14",2007,4.6,"Tübingen"
"Y_GE15","DE2",2007,5.3,"Bayern"
"Y_GE15","DE21",2007,4.4,"Oberbayern"
"Y_GE15","DE22",2007,5,"Niederbayern"
"Y_GE15","DE23",2007,5.3,"Oberpfalz"
"Y_GE15","DE24",2007,7.7,"Oberfranken"
"Y_GE15","DE25",2007,6.7,"Mittelfranken"
"Y_GE15","DE26",2007,5.8,"Unterfranken"
"Y_GE15","DE27",2007,5,"Schwaben"
"Y_GE15","DE3",2007,16.4,"Berlin"
"Y_GE15","DE30",2007,16.4,"Berlin"
"Y_GE15","DE4",2007,13.8,"Brandenburg"
"Y_GE15","DE40",2007,13.8,"Brandenburg"
"Y_GE15","DE5",2007,11.9,"Bremen"
"Y_GE15","DE50",2007,11.9,"Bremen"
"Y_GE15","DE6",2007,9,"Hamburg"
"Y_GE15","DE60",2007,9,"Hamburg"
"Y_GE15","DE7",2007,7.3,"Hessen"
"Y_GE15","DE71",2007,7.2,"Darmstadt"
"Y_GE15","DE72",2007,7.2,"Gießen"
"Y_GE15","DE73",2007,8,"Kassel"
"Y_GE15","DE8",2007,17.5,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2007,17.5,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2007,7.9,"Niedersachsen"
"Y_GE15","DE91",2007,8.9,"Braunschweig"
"Y_GE15","DE92",2007,8.4,"Hannover"
"Y_GE15","DE93",2007,7.4,"Lüneburg"
"Y_GE15","DE94",2007,7.1,"Weser-Ems"
"Y_GE15","DEA",2007,8.4,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2007,8.6,"Düsseldorf"
"Y_GE15","DEA2",2007,7.7,"Köln"
"Y_GE15","DEA3",2007,7.3,"Münster"
"Y_GE15","DEA4",2007,8.1,"Detmold"
"Y_GE15","DEA5",2007,9.7,"Arnsberg"
"Y_GE15","DEB",2007,6,"Rheinland-Pfalz"
"Y_GE15","DEB1",2007,6.3,"Koblenz"
"Y_GE15","DEB2",2007,5.3,"Trier"
"Y_GE15","DEB3",2007,5.9,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2007,7.3,"Saarland"
"Y_GE15","DEC0",2007,7.3,"Saarland"
"Y_GE15","DED",2007,14.5,"Sachsen"
"Y_GE15","DED2",2007,13.4,"Dresden"
"Y_GE15","DED4",2007,13.9,"Chemnitz"
"Y_GE15","DED5",2007,17.3,"Leipzig"
"Y_GE15","DEE",2007,15.7,"Sachsen-Anhalt"
"Y_GE15","DEE0",2007,15.7,"Sachsen-Anhalt"
"Y_GE15","DEF",2007,8,"Schleswig-Holstein"
"Y_GE15","DEF0",2007,8,"Schleswig-Holstein"
"Y_GE15","DEG",2007,13.8,"Thüringen"
"Y_GE15","DEG0",2007,13.8,"Thüringen"
"Y_GE15","DK",2007,3.8,"Denmark"
"Y_GE15","DK0",2007,3.8,"Danmark"
"Y_GE15","DK01",2007,4.3,"Hovedstaden"
"Y_GE15","DK02",2007,3.6,"Sjælland"
"Y_GE15","DK03",2007,3.5,"Syddanmark"
"Y_GE15","DK04",2007,3.3,"Midtjylland"
"Y_GE15","DK05",2007,4.4,"Nordjylland"
"Y_GE15","EA17",2007,7.5,"Euro area (17 countries)"
"Y_GE15","EA18",2007,7.5,"Euro area (18 countries)"
"Y_GE15","EA19",2007,7.4,"Euro area (19 countries)"
"Y_GE15","EE",2007,4.6,"Estonia"
"Y_GE15","EE0",2007,4.6,"Eesti"
"Y_GE15","EE00",2007,4.6,"Eesti"
"Y_GE15","EL",2007,8.4,"Greece"
"Y_GE15","EL1",2007,9.2,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2007,9.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2007,9.1,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2007,12.1,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2007,7.8,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2007,9.1,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2007,10,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2007,9,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2007,9.9,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2007,9.4,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2007,7.3,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2007,7.8,"Attiki"
"Y_GE15","EL30",2007,7.8,"Attiki"
"Y_GE15","EL4",2007,7,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2007,8.1,"Voreio Aigaio"
"Y_GE15","EL42",2007,9.4,"Notio Aigaio"
"Y_GE15","EL43",2007,5.4,"Kriti"
"Y_GE15","ES",2007,8.2,"Spain"
"Y_GE15","ES1",2007,7.5,"Noroeste (ES)"
"Y_GE15","ES11",2007,7.6,"Galicia"
"Y_GE15","ES12",2007,8.4,"Principado de Asturias"
"Y_GE15","ES13",2007,6,"Cantabria"
"Y_GE15","ES2",2007,5.7,"Noreste (ES)"
"Y_GE15","ES21",2007,6.2,"País Vasco"
"Y_GE15","ES22",2007,4.7,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2007,5.8,"La Rioja"
"Y_GE15","ES24",2007,5.3,"Aragón"
"Y_GE15","ES3",2007,6.2,"Comunidad de Madrid"
"Y_GE15","ES30",2007,6.2,"Comunidad de Madrid"
"Y_GE15","ES4",2007,8.4,"Centro (ES)"
"Y_GE15","ES41",2007,7.1,"Castilla y León"
"Y_GE15","ES42",2007,7.7,"Castilla-la Mancha"
"Y_GE15","ES43",2007,13,"Extremadura"
"Y_GE15","ES5",2007,7.3,"Este (ES)"
"Y_GE15","ES51",2007,6.5,"Cataluña"
"Y_GE15","ES52",2007,8.7,"Comunidad Valenciana"
"Y_GE15","ES53",2007,7.2,"Illes Balears"
"Y_GE15","ES6",2007,12,"Sur (ES)"
"Y_GE15","ES61",2007,12.8,"Andalucía"
"Y_GE15","ES62",2007,7.5,"Región de Murcia"
"Y_GE15","ES63",2007,21,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2007,18.2,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2007,10.5,"Canarias (ES)"
"Y_GE15","ES70",2007,10.5,"Canarias (ES)"
"Y_GE15","EU15",2007,7,"European Union (15 countries)"
"Y_GE15","EU27",2007,7.1,"European Union (27 countries)"
"Y_GE15","EU28",2007,7.2,"European Union (28 countries)"
"Y_GE15","FI",2007,6.9,"Finland"
"Y_GE15","FI1",2007,6.9,"Manner-Suomi"
"Y_GE15","FI19",2007,6.5,"Länsi-Suomi"
"Y_GE15","FI1B",2007,5,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2007,6.7,"Etelä-Suomi"
"Y_GE15","FI1D",2007,9.9,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2007,NA,"Åland"
"Y_GE15","FI20",2007,NA,"Åland"
"Y_GE15","FR",2007,8,"France"
"Y_GE15","FR1",2007,7.8,"Île de France"
"Y_GE15","FR10",2007,7.8,"Île de France"
"Y_GE15","FR2",2007,7.4,"Bassin Parisien"
"Y_GE15","FR21",2007,8,"Champagne-Ardenne"
"Y_GE15","FR22",2007,9.9,"Picardie"
"Y_GE15","FR23",2007,8.6,"Haute-Normandie"
"Y_GE15","FR24",2007,5.8,"Centre (FR)"
"Y_GE15","FR25",2007,5.6,"Basse-Normandie"
"Y_GE15","FR26",2007,6.7,"Bourgogne"
"Y_GE15","FR3",2007,11.3,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2007,11.3,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2007,6.8,"Est (FR)"
"Y_GE15","FR41",2007,7.5,"Lorraine"
"Y_GE15","FR42",2007,5.9,"Alsace"
"Y_GE15","FR43",2007,7.1,"Franche-Comté"
"Y_GE15","FR5",2007,6.3,"Ouest (FR)"
"Y_GE15","FR51",2007,5.9,"Pays de la Loire"
"Y_GE15","FR52",2007,6.7,"Bretagne"
"Y_GE15","FR53",2007,6.5,"Poitou-Charentes"
"Y_GE15","FR6",2007,7.3,"Sud-Ouest (FR)"
"Y_GE15","FR61",2007,6.9,"Aquitaine"
"Y_GE15","FR62",2007,7.9,"Midi-Pyrénées"
"Y_GE15","FR63",2007,6.7,"Limousin"
"Y_GE15","FR7",2007,6.7,"Centre-Est (FR)"
"Y_GE15","FR71",2007,6.3,"Rhône-Alpes"
"Y_GE15","FR72",2007,8.3,"Auvergne"
"Y_GE15","FR8",2007,9.4,"Méditerranée"
"Y_GE15","FR81",2007,10.1,"Languedoc-Roussillon"
"Y_GE15","FR82",2007,9,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2007,11.1,"Corse"
"Y_GE15","FR9",2007,22.7,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2007,22.6,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2007,21.1,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2007,20.1,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2007,24.1,"Réunion (NUTS 2010)"
"Y_GE15","HR",2007,9.9,"Croatia"
"Y_GE15","HR0",2007,9.9,"Hrvatska"
"Y_GE15","HR03",2007,9.2,"Jadranska Hrvatska"
"Y_GE15","HR04",2007,10.3,"Kontinentalna Hrvatska"
"Y_GE15","HU",2007,7.4,"Hungary"
"Y_GE15","HU1",2007,4.8,"Közép-Magyarország"
"Y_GE15","HU10",2007,4.8,"Közép-Magyarország"
"Y_GE15","HU2",2007,6.4,"Dunántúl"
"Y_GE15","HU21",2007,4.9,"Közép-Dunántúl"
"Y_GE15","HU22",2007,5.1,"Nyugat-Dunántúl"
"Y_GE15","HU23",2007,9.9,"Dél-Dunántúl"
"Y_GE15","HU3",2007,10.4,"Alföld és Észak"
"Y_GE15","HU31",2007,12.6,"Észak-Magyarország"
"Y_GE15","HU32",2007,10.7,"Észak-Alföld"
"Y_GE15","HU33",2007,8,"Dél-Alföld"
"Y_GE15","IE",2007,4.7,"Ireland"
"Y_GE15","IE0",2007,4.7,"Éire/Ireland"
"Y_GE15","IE01",2007,5,"Border, Midland and Western"
"Y_GE15","IE02",2007,4.6,"Southern and Eastern"
"Y_GE15","IS",2007,2.3,"Iceland"
"Y_GE15","IS0",2007,2.3,"Ísland"
"Y_GE15","IS00",2007,2.3,"Ísland"
"Y_GE15","IT",2007,6.1,"Italy"
"Y_GE15","ITC",2007,3.8,"Nord-Ovest"
"Y_GE15","ITC1",2007,4.2,"Piemonte"
"Y_GE15","ITC2",2007,3.2,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2007,4.8,"Liguria"
"Y_GE15","ITC4",2007,3.4,"Lombardia"
"Y_GE15","ITF",2007,10.4,"Sud"
"Y_GE15","ITF1",2007,6.2,"Abruzzo"
"Y_GE15","ITF2",2007,8.1,"Molise"
"Y_GE15","ITF3",2007,11.2,"Campania"
"Y_GE15","ITF4",2007,11.1,"Puglia"
"Y_GE15","ITF5",2007,9.4,"Basilicata"
"Y_GE15","ITF6",2007,11.1,"Calabria"
"Y_GE15","ITG",2007,12,"Isole"
"Y_GE15","ITG1",2007,12.9,"Sicilia"
"Y_GE15","ITG2",2007,9.8,"Sardegna"
"Y_GE15","ITH",2007,3.1,"Nord-Est"
"Y_GE15","ITH1",2007,2.6,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2007,2.9,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2007,3.4,"Veneto"
"Y_GE15","ITH4",2007,3.4,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2007,2.8,"Emilia-Romagna"
"Y_GE15","ITI",2007,5.3,"Centro (IT)"
"Y_GE15","ITI1",2007,4.4,"Toscana"
"Y_GE15","ITI2",2007,4.6,"Umbria"
"Y_GE15","ITI3",2007,4.1,"Marche"
"Y_GE15","ITI4",2007,6.4,"Lazio"
"Y_GE15","LT",2007,4.2,"Lithuania"
"Y_GE15","LT0",2007,4.2,"Lietuva"
"Y_GE15","LT00",2007,4.2,"Lietuva"
"Y_GE15","LU",2007,4.1,"Luxembourg"
"Y_GE15","LU0",2007,4.1,"Luxembourg"
"Y_GE15","LU00",2007,4.1,"Luxembourg"
"Y_GE15","LV",2007,6.1,"Latvia"
"Y_GE15","LV0",2007,6.1,"Latvija"
"Y_GE15","LV00",2007,6.1,"Latvija"
"Y_GE15","MK",2007,34.9,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2007,34.9,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2007,34.9,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2007,6.5,"Malta"
"Y_GE15","MT0",2007,6.5,"Malta"
"Y_GE15","MT00",2007,6.5,"Malta"
"Y_GE15","NL",2007,3.2,"Netherlands"
"Y_GE15","NL1",2007,3.9,"Noord-Nederland"
"Y_GE15","NL11",2007,4.9,"Groningen"
"Y_GE15","NL12",2007,3.2,"Friesland (NL)"
"Y_GE15","NL13",2007,3.7,"Drenthe"
"Y_GE15","NL2",2007,3,"Oost-Nederland"
"Y_GE15","NL21",2007,3.2,"Overijssel"
"Y_GE15","NL22",2007,2.7,"Gelderland"
"Y_GE15","NL23",2007,4.1,"Flevoland"
"Y_GE15","NL3",2007,3.1,"West-Nederland"
"Y_GE15","NL31",2007,2.7,"Utrecht"
"Y_GE15","NL32",2007,2.9,"Noord-Holland"
"Y_GE15","NL33",2007,3.5,"Zuid-Holland"
"Y_GE15","NL34",2007,2.1,"Zeeland"
"Y_GE15","NL4",2007,3.1,"Zuid-Nederland"
"Y_GE15","NL41",2007,2.8,"Noord-Brabant"
"Y_GE15","NL42",2007,3.9,"Limburg (NL)"
"Y_GE15","NO",2007,2.5,"Norway"
"Y_GE15","NO0",2007,2.5,"Norge"
"Y_GE15","NO01",2007,2.5,"Oslo og Akershus"
"Y_GE15","NO02",2007,2.2,"Hedmark og Oppland"
"Y_GE15","NO03",2007,2.9,"Sør-Østlandet"
"Y_GE15","NO04",2007,1.9,"Agder og Rogaland"
"Y_GE15","NO05",2007,2.3,"Vestlandet"
"Y_GE15","NO06",2007,3.1,"Trøndelag"
"Y_GE15","NO07",2007,2.7,"Nord-Norge"
"Y_GE15","PL",2007,9.6,"Poland"
"Y_GE15","PL1",2007,9.1,"Region Centralny"
"Y_GE15","PL11",2007,9.3,"Lódzkie"
"Y_GE15","PL12",2007,9.1,"Mazowieckie"
"Y_GE15","PL2",2007,8.3,"Region Poludniowy"
"Y_GE15","PL21",2007,8.5,"Malopolskie"
"Y_GE15","PL22",2007,8.1,"Slaskie"
"Y_GE15","PL3",2007,10,"Region Wschodni"
"Y_GE15","PL31",2007,9.5,"Lubelskie"
"Y_GE15","PL32",2007,9.6,"Podkarpackie"
"Y_GE15","PL33",2007,12.1,"Swietokrzyskie"
"Y_GE15","PL34",2007,8.9,"Podlaskie"
"Y_GE15","PL4",2007,9.3,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2007,8.3,"Wielkopolskie"
"Y_GE15","PL42",2007,11.5,"Zachodniopomorskie"
"Y_GE15","PL43",2007,9.8,"Lubuskie"
"Y_GE15","PL5",2007,11.9,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2007,12.7,"Dolnoslaskie"
"Y_GE15","PL52",2007,9.4,"Opolskie"
"Y_GE15","PL6",2007,10.4,"Region Pólnocny"
"Y_GE15","PL61",2007,11.3,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2007,10.5,"Warminsko-Mazurskie"
"Y_GE15","PL63",2007,9.5,"Pomorskie"
"Y_GE15","PT",2007,8,"Portugal"
"Y_GE15","PT1",2007,8.1,"Continente"
"Y_GE15","PT11",2007,9.3,"Norte"
"Y_GE15","PT15",2007,6.7,"Algarve"
"Y_GE15","PT16",2007,5.5,"Centro (PT)"
"Y_GE15","PT17",2007,8.9,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2007,8.4,"Alentejo"
"Y_GE15","PT2",2007,4.3,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2007,4.3,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2007,6.8,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2007,6.8,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2007,6.4,"Romania"
"Y_GE15","RO1",2007,6.3,"Macroregiunea unu"
"Y_GE15","RO11",2007,4.3,"Nord-Vest"
"Y_GE15","RO12",2007,8.5,"Centru"
"Y_GE15","RO2",2007,6.5,"Macroregiunea doi"
"Y_GE15","RO21",2007,5,"Nord-Est"
"Y_GE15","RO22",2007,8.5,"Sud-Est"
"Y_GE15","RO3",2007,6.6,"Macroregiunea trei"
"Y_GE15","RO31",2007,8.2,"Sud - Muntenia"
"Y_GE15","RO32",2007,4.1,"Bucuresti - Ilfov"
"Y_GE15","RO4",2007,6.3,"Macroregiunea patru"
"Y_GE15","RO41",2007,6.8,"Sud-Vest Oltenia"
"Y_GE15","RO42",2007,5.6,"Vest"
"Y_GE15","SE",2007,6.2,"Sweden"
"Y_GE15","SE1",2007,6.1,"Östra Sverige"
"Y_GE15","SE11",2007,5.6,"Stockholm"
"Y_GE15","SE12",2007,6.7,"Östra Mellansverige"
"Y_GE15","SE2",2007,6.1,"Södra Sverige"
"Y_GE15","SE21",2007,5.1,"Småland med öarna"
"Y_GE15","SE22",2007,7.1,"Sydsverige"
"Y_GE15","SE23",2007,5.9,"Västsverige"
"Y_GE15","SE3",2007,6.5,"Norra Sverige"
"Y_GE15","SE31",2007,6.3,"Norra Mellansverige"
"Y_GE15","SE32",2007,6.3,"Mellersta Norrland"
"Y_GE15","SE33",2007,6.8,"Övre Norrland"
"Y_GE15","SI",2007,4.8,"Slovenia"
"Y_GE15","SI0",2007,4.8,"Slovenija"
"Y_GE15","SI01",2007,5.6,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2007,3.9,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2007,11.1,"Slovakia"
"Y_GE15","SK0",2007,11.1,"Slovensko"
"Y_GE15","SK01",2007,4.3,"Bratislavský kraj"
"Y_GE15","SK02",2007,7.8,"Západné Slovensko"
"Y_GE15","SK03",2007,15.3,"Stredné Slovensko"
"Y_GE15","SK04",2007,14.9,"Východné Slovensko"
"Y_GE15","TR",2007,8.9,"Turkey"
"Y_GE15","TR1",2007,9.4,"Istanbul"
"Y_GE15","TR10",2007,9.4,"Istanbul"
"Y_GE15","TR2",2007,5.5,"Bati Marmara"
"Y_GE15","TR21",2007,6.5,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2007,4.6,"Balikesir, Çanakkale"
"Y_GE15","TR3",2007,7.9,"Ege"
"Y_GE15","TR31",2007,9.3,"Izmir"
"Y_GE15","TR32",2007,8.2,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2007,5.6,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2007,8.6,"Dogu Marmara"
"Y_GE15","TR41",2007,7.4,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2007,10.2,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2007,10,"Bati Anadolu"
"Y_GE15","TR51",2007,10.5,"Ankara"
"Y_GE15","TR52",2007,8.9,"Konya, Karaman"
"Y_GE15","TR6",2007,9.9,"Akdeniz"
"Y_GE15","TR61",2007,6.2,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2007,13,"Adana, Mersin"
"Y_GE15","TR63",2007,9.7,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2007,8.8,"Orta Anadolu"
"Y_GE15","TR71",2007,7.1,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2007,9.9,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2007,6.5,"Bati Karadeniz"
"Y_GE15","TR81",2007,7,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2007,3.2,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2007,7.1,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2007,4.9,"Dogu Karadeniz"
"Y_GE15","TR90",2007,4.9,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2007,4.3,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2007,4.3,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2007,4.4,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2007,11,"Ortadogu Anadolu"
"Y_GE15","TRB1",2007,10.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2007,11.4,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2007,15.7,"Güneydogu Anadolu"
"Y_GE15","TRC1",2007,16.9,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2007,12.9,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2007,18,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2007,5.3,"United Kingdom"
"Y_GE15","UKC",2007,6.1,"North East (UK)"
"Y_GE15","UKC1",2007,6,"Tees Valley and Durham"
"Y_GE15","UKC2",2007,6.2,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2007,5.8,"North West (UK)"
"Y_GE15","UKD1",2007,3.3,"Cumbria"
"Y_GE15","UKD3",2007,6.4,"Greater Manchester"
"Y_GE15","UKD4",2007,5.6,"Lancashire"
"Y_GE15","UKD6",2007,2.9,"Cheshire"
"Y_GE15","UKD7",2007,7.6,"Merseyside"
"Y_GE15","UKE",2007,5.5,"Yorkshire and The Humber"
"Y_GE15","UKE1",2007,6.1,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2007,3.4,"North Yorkshire"
"Y_GE15","UKE3",2007,6.2,"South Yorkshire"
"Y_GE15","UKE4",2007,5.6,"West Yorkshire"
"Y_GE15","UKF",2007,5.2,"East Midlands (UK)"
"Y_GE15","UKF1",2007,5.8,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2007,4.6,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2007,5.4,"Lincolnshire"
"Y_GE15","UKG",2007,6.2,"West Midlands (UK)"
"Y_GE15","UKG1",2007,3.9,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2007,5.3,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2007,8.1,"West Midlands"
"Y_GE15","UKH",2007,4.6,"East of England"
"Y_GE15","UKH1",2007,4.3,"East Anglia"
"Y_GE15","UKH2",2007,4.7,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2007,5,"Essex"
"Y_GE15","UKI",2007,6.8,"London"
"Y_GE15","UKI1",2007,8.2,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2007,5.9,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2007,4.4,"South East (UK)"
"Y_GE15","UKJ1",2007,4,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2007,4,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2007,4.3,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2007,5.6,"Kent"
"Y_GE15","UKK",2007,3.8,"South West (UK)"
"Y_GE15","UKK1",2007,3.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2007,3.7,"Dorset and Somerset"
"Y_GE15","UKK3",2007,4.4,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2007,4.7,"Devon"
"Y_GE15","UKL",2007,5.2,"Wales"
"Y_GE15","UKL1",2007,5.5,"West Wales and The Valleys"
"Y_GE15","UKL2",2007,4.8,"East Wales"
"Y_GE15","UKM",2007,4.7,"Scotland"
"Y_GE15","UKM2",2007,5.1,"Eastern Scotland"
"Y_GE15","UKM3",2007,5.2,"South Western Scotland"
"Y_GE15","UKM5",2007,3.3,"North Eastern Scotland"
"Y_GE15","UKM6",2007,2.2,"Highlands and Islands"
"Y_GE15","UKN",2007,3.8,"Northern Ireland (UK)"
"Y_GE15","UKN0",2007,3.8,"Northern Ireland (UK)"
"Y_GE25","AT",2007,4.1,"Austria"
"Y_GE25","AT1",2007,5.6,"Ostösterreich"
"Y_GE25","AT11",2007,3.4,"Burgenland (AT)"
"Y_GE25","AT12",2007,3.3,"Niederösterreich"
"Y_GE25","AT13",2007,8.1,"Wien"
"Y_GE25","AT2",2007,3.4,"Südösterreich"
"Y_GE25","AT21",2007,3.5,"Kärnten"
"Y_GE25","AT22",2007,3.3,"Steiermark"
"Y_GE25","AT3",2007,2.8,"Westösterreich"
"Y_GE25","AT31",2007,2.8,"Oberösterreich"
"Y_GE25","AT32",2007,3.1,"Salzburg"
"Y_GE25","AT33",2007,2.3,"Tirol"
"Y_GE25","AT34",2007,3.2,"Vorarlberg"
"Y_GE25","BE",2007,6.3,"Belgium"
"Y_GE25","BE1",2007,15.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2007,15.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2007,3.6,"Vlaams Gewest"
"Y_GE25","BE21",2007,4.4,"Prov. Antwerpen"
"Y_GE25","BE22",2007,4.5,"Prov. Limburg (BE)"
"Y_GE25","BE23",2007,3.9,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2007,2.6,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2007,2.3,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2007,8.6,"Région wallonne"
"Y_GE25","BE31",2007,6,"Prov. Brabant Wallon"
"Y_GE25","BE32",2007,10.3,"Prov. Hainaut"
"Y_GE25","BE33",2007,9.3,"Prov. Liège"
"Y_GE25","BE34",2007,5.5,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2007,6.8,"Prov. Namur"
"Y_GE25","BG",2007,6.1,"Bulgaria"
"Y_GE25","BG3",2007,8.1,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2007,7.9,"Severozapaden"
"Y_GE25","BG32",2007,9.7,"Severen tsentralen"
"Y_GE25","BG33",2007,9.4,"Severoiztochen"
"Y_GE25","BG34",2007,5.8,"Yugoiztochen"
"Y_GE25","BG4",2007,4.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2007,3.7,"Yugozapaden"
"Y_GE25","BG42",2007,4.9,"Yuzhen tsentralen"
"Y_GE25","CH",2007,3.1,"Switzerland"
"Y_GE25","CH0",2007,3.1,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2007,4.1,"Région lémanique"
"Y_GE25","CH02",2007,3.2,"Espace Mittelland"
"Y_GE25","CH03",2007,2.7,"Nordwestschweiz"
"Y_GE25","CH04",2007,2.9,"Zürich"
"Y_GE25","CH05",2007,2.3,"Ostschweiz"
"Y_GE25","CH06",2007,2.4,"Zentralschweiz"
"Y_GE25","CH07",2007,4.3,"Ticino"
"Y_GE25","CY",2007,3.2,"Cyprus"
"Y_GE25","CY0",2007,3.2,"Kypros"
"Y_GE25","CY00",2007,3.2,"Kypros"
"Y_GE25","CZ",2007,4.8,"Czech Republic"
"Y_GE25","CZ0",2007,4.8,"Ceská republika"
"Y_GE25","CZ01",2007,2.2,"Praha"
"Y_GE25","CZ02",2007,3,"Strední Cechy"
"Y_GE25","CZ03",2007,3.3,"Jihozápad"
"Y_GE25","CZ04",2007,8.4,"Severozápad"
"Y_GE25","CZ05",2007,4.4,"Severovýchod"
"Y_GE25","CZ06",2007,4.6,"Jihovýchod"
"Y_GE25","CZ07",2007,5.7,"Strední Morava"
"Y_GE25","CZ08",2007,7.9,"Moravskoslezsko"
"Y_GE25","DE",2007,8.2,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2007,4.7,"Baden-Württemberg"
"Y_GE25","DE11",2007,4.7,"Stuttgart"
"Y_GE25","DE12",2007,5.3,"Karlsruhe"
"Y_GE25","DE13",2007,4.2,"Freiburg"
"Y_GE25","DE14",2007,4.3,"Tübingen"
"Y_GE25","DE2",2007,5,"Bayern"
"Y_GE25","DE21",2007,4.1,"Oberbayern"
"Y_GE25","DE22",2007,4.7,"Niederbayern"
"Y_GE25","DE23",2007,4.9,"Oberpfalz"
"Y_GE25","DE24",2007,7.1,"Oberfranken"
"Y_GE25","DE25",2007,6.3,"Mittelfranken"
"Y_GE25","DE26",2007,5.1,"Unterfranken"
"Y_GE25","DE27",2007,4.8,"Schwaben"
"Y_GE25","DE3",2007,15.8,"Berlin"
"Y_GE25","DE30",2007,15.8,"Berlin"
"Y_GE25","DE4",2007,13.4,"Brandenburg"
"Y_GE25","DE40",2007,13.4,"Brandenburg"
"Y_GE25","DE5",2007,12.2,"Bremen"
"Y_GE25","DE50",2007,12.2,"Bremen"
"Y_GE25","DE6",2007,8.7,"Hamburg"
"Y_GE25","DE60",2007,8.7,"Hamburg"
"Y_GE25","DE7",2007,6.8,"Hessen"
"Y_GE25","DE71",2007,6.7,"Darmstadt"
"Y_GE25","DE72",2007,6.3,"Gießen"
"Y_GE25","DE73",2007,7.3,"Kassel"
"Y_GE25","DE8",2007,17.1,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2007,17.1,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2007,7.4,"Niedersachsen"
"Y_GE25","DE91",2007,8.4,"Braunschweig"
"Y_GE25","DE92",2007,7.8,"Hannover"
"Y_GE25","DE93",2007,7,"Lüneburg"
"Y_GE25","DE94",2007,6.6,"Weser-Ems"
"Y_GE25","DEA",2007,7.8,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2007,7.9,"Düsseldorf"
"Y_GE25","DEA2",2007,7.3,"Köln"
"Y_GE25","DEA3",2007,7.1,"Münster"
"Y_GE25","DEA4",2007,7.6,"Detmold"
"Y_GE25","DEA5",2007,9.1,"Arnsberg"
"Y_GE25","DEB",2007,5.3,"Rheinland-Pfalz"
"Y_GE25","DEB1",2007,5.8,"Koblenz"
"Y_GE25","DEB2",2007,4.8,"Trier"
"Y_GE25","DEB3",2007,5.1,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2007,7.1,"Saarland"
"Y_GE25","DEC0",2007,7.1,"Saarland"
"Y_GE25","DED",2007,14.3,"Sachsen"
"Y_GE25","DED2",2007,13,"Dresden"
"Y_GE25","DED4",2007,13.8,"Chemnitz"
"Y_GE25","DED5",2007,17.1,"Leipzig"
"Y_GE25","DEE",2007,15.1,"Sachsen-Anhalt"
"Y_GE25","DEE0",2007,15.1,"Sachsen-Anhalt"
"Y_GE25","DEF",2007,7.3,"Schleswig-Holstein"
"Y_GE25","DEF0",2007,7.3,"Schleswig-Holstein"
"Y_GE25","DEG",2007,13.6,"Thüringen"
"Y_GE25","DEG0",2007,13.6,"Thüringen"
"Y_GE25","DK",2007,3.2,"Denmark"
"Y_GE25","DK0",2007,3.2,"Danmark"
"Y_GE25","DK01",2007,3.8,"Hovedstaden"
"Y_GE25","DK02",2007,2.9,"Sjælland"
"Y_GE25","DK03",2007,2.7,"Syddanmark"
"Y_GE25","DK04",2007,2.7,"Midtjylland"
"Y_GE25","DK05",2007,3.5,"Nordjylland"
"Y_GE25","EA17",2007,6.5,"Euro area (17 countries)"
"Y_GE25","EA18",2007,6.5,"Euro area (18 countries)"
"Y_GE25","EA19",2007,6.5,"Euro area (19 countries)"
"Y_GE25","EE",2007,3.9,"Estonia"
"Y_GE25","EE0",2007,3.9,"Eesti"
"Y_GE25","EE00",2007,3.9,"Eesti"
"Y_GE25","EL",2007,7.2,"Greece"
"Y_GE25","EL1",2007,7.9,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2007,8.2,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2007,7.9,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2007,10.7,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2007,6.5,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2007,7.5,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2007,8.5,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2007,7.7,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2007,7.8,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2007,7.8,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2007,6.1,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2007,6.7,"Attiki"
"Y_GE25","EL30",2007,6.7,"Attiki"
"Y_GE25","EL4",2007,6,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2007,5.6,"Voreio Aigaio"
"Y_GE25","EL42",2007,9,"Notio Aigaio"
"Y_GE25","EL43",2007,4.7,"Kriti"
"Y_GE25","ES",2007,7,"Spain"
"Y_GE25","ES1",2007,6.7,"Noroeste (ES)"
"Y_GE25","ES11",2007,6.8,"Galicia"
"Y_GE25","ES12",2007,7.5,"Principado de Asturias"
"Y_GE25","ES13",2007,5.2,"Cantabria"
"Y_GE25","ES2",2007,4.8,"Noreste (ES)"
"Y_GE25","ES21",2007,5.3,"País Vasco"
"Y_GE25","ES22",2007,4,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2007,4.5,"La Rioja"
"Y_GE25","ES24",2007,4.4,"Aragón"
"Y_GE25","ES3",2007,5,"Comunidad de Madrid"
"Y_GE25","ES30",2007,5,"Comunidad de Madrid"
"Y_GE25","ES4",2007,7.1,"Centro (ES)"
"Y_GE25","ES41",2007,6.1,"Castilla y León"
"Y_GE25","ES42",2007,6.4,"Castilla-la Mancha"
"Y_GE25","ES43",2007,11.1,"Extremadura"
"Y_GE25","ES5",2007,6.3,"Este (ES)"
"Y_GE25","ES51",2007,5.7,"Cataluña"
"Y_GE25","ES52",2007,7.4,"Comunidad Valenciana"
"Y_GE25","ES53",2007,6.2,"Illes Balears"
"Y_GE25","ES6",2007,10.5,"Sur (ES)"
"Y_GE25","ES61",2007,11.1,"Andalucía"
"Y_GE25","ES62",2007,6.2,"Región de Murcia"
"Y_GE25","ES63",2007,18.1,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2007,16.1,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2007,9,"Canarias (ES)"
"Y_GE25","ES70",2007,9,"Canarias (ES)"
"Y_GE25","EU15",2007,6,"European Union (15 countries)"
"Y_GE25","EU27",2007,6.1,"European Union (27 countries)"
"Y_GE25","EU28",2007,6.1,"European Union (28 countries)"
"Y_GE25","FI",2007,5.4,"Finland"
"Y_GE25","FI1",2007,5.5,"Manner-Suomi"
"Y_GE25","FI19",2007,5.2,"Länsi-Suomi"
"Y_GE25","FI1B",2007,3.9,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2007,5.4,"Etelä-Suomi"
"Y_GE25","FI1D",2007,7.9,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2007,NA,"Åland"
"Y_GE25","FI20",2007,NA,"Åland"
"Y_GE25","FR",2007,6.7,"France"
"Y_GE25","FR1",2007,6.7,"Île de France"
"Y_GE25","FR10",2007,6.7,"Île de France"
"Y_GE25","FR2",2007,5.9,"Bassin Parisien"
"Y_GE25","FR21",2007,6.1,"Champagne-Ardenne"
"Y_GE25","FR22",2007,8.1,"Picardie"
"Y_GE25","FR23",2007,6.3,"Haute-Normandie"
"Y_GE25","FR24",2007,4.9,"Centre (FR)"
"Y_GE25","FR25",2007,4.5,"Basse-Normandie"
"Y_GE25","FR26",2007,5.7,"Bourgogne"
"Y_GE25","FR3",2007,9,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2007,9,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2007,5.5,"Est (FR)"
"Y_GE25","FR41",2007,6.2,"Lorraine"
"Y_GE25","FR42",2007,4.6,"Alsace"
"Y_GE25","FR43",2007,5.9,"Franche-Comté"
"Y_GE25","FR5",2007,5.5,"Ouest (FR)"
"Y_GE25","FR51",2007,5.2,"Pays de la Loire"
"Y_GE25","FR52",2007,5.9,"Bretagne"
"Y_GE25","FR53",2007,5.2,"Poitou-Charentes"
"Y_GE25","FR6",2007,5.9,"Sud-Ouest (FR)"
"Y_GE25","FR61",2007,5.5,"Aquitaine"
"Y_GE25","FR62",2007,6.4,"Midi-Pyrénées"
"Y_GE25","FR63",2007,5.6,"Limousin"
"Y_GE25","FR7",2007,5.4,"Centre-Est (FR)"
"Y_GE25","FR71",2007,5.2,"Rhône-Alpes"
"Y_GE25","FR72",2007,6.8,"Auvergne"
"Y_GE25","FR8",2007,8,"Méditerranée"
"Y_GE25","FR81",2007,8.5,"Languedoc-Roussillon"
"Y_GE25","FR82",2007,7.7,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2007,9.3,"Corse"
"Y_GE25","FR9",2007,19.8,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2007,20.2,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2007,19.1,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2007,17.9,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2007,20.4,"Réunion (NUTS 2010)"
"Y_GE25","HR",2007,8.2,"Croatia"
"Y_GE25","HR0",2007,8.2,"Hrvatska"
"Y_GE25","HR03",2007,7.9,"Jadranska Hrvatska"
"Y_GE25","HR04",2007,8.4,"Kontinentalna Hrvatska"
"Y_GE25","HU",2007,6.5,"Hungary"
"Y_GE25","HU1",2007,4.4,"Közép-Magyarország"
"Y_GE25","HU10",2007,4.4,"Közép-Magyarország"
"Y_GE25","HU2",2007,5.7,"Dunántúl"
"Y_GE25","HU21",2007,4.3,"Közép-Dunántúl"
"Y_GE25","HU22",2007,4.5,"Nyugat-Dunántúl"
"Y_GE25","HU23",2007,8.8,"Dél-Dunántúl"
"Y_GE25","HU3",2007,9,"Alföld és Észak"
"Y_GE25","HU31",2007,11.1,"Észak-Magyarország"
"Y_GE25","HU32",2007,9.2,"Észak-Alföld"
"Y_GE25","HU33",2007,7.1,"Dél-Alföld"
"Y_GE25","IE",2007,3.8,"Ireland"
"Y_GE25","IE0",2007,3.8,"Éire/Ireland"
"Y_GE25","IE01",2007,4,"Border, Midland and Western"
"Y_GE25","IE02",2007,3.7,"Southern and Eastern"
"Y_GE25","IS",2007,1.3,"Iceland"
"Y_GE25","IS0",2007,1.3,"Ísland"
"Y_GE25","IS00",2007,1.3,"Ísland"
"Y_GE25","IT",2007,4.9,"Italy"
"Y_GE25","ITC",2007,3,"Nord-Ovest"
"Y_GE25","ITC1",2007,3.5,"Piemonte"
"Y_GE25","ITC2",2007,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2007,3.9,"Liguria"
"Y_GE25","ITC4",2007,2.7,"Lombardia"
"Y_GE25","ITF",2007,8.5,"Sud"
"Y_GE25","ITF1",2007,5.3,"Abruzzo"
"Y_GE25","ITF2",2007,6.7,"Molise"
"Y_GE25","ITF3",2007,9,"Campania"
"Y_GE25","ITF4",2007,8.7,"Puglia"
"Y_GE25","ITF5",2007,7.7,"Basilicata"
"Y_GE25","ITF6",2007,9.4,"Calabria"
"Y_GE25","ITG",2007,9.6,"Isole"
"Y_GE25","ITG1",2007,10.4,"Sicilia"
"Y_GE25","ITG2",2007,7.8,"Sardegna"
"Y_GE25","ITH",2007,2.6,"Nord-Est"
"Y_GE25","ITH1",2007,2.2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2007,2.4,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2007,3,"Veneto"
"Y_GE25","ITH4",2007,2.6,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2007,2.3,"Emilia-Romagna"
"Y_GE25","ITI",2007,4.4,"Centro (IT)"
"Y_GE25","ITI1",2007,3.7,"Toscana"
"Y_GE25","ITI2",2007,4,"Umbria"
"Y_GE25","ITI3",2007,3.7,"Marche"
"Y_GE25","ITI4",2007,5.1,"Lazio"
"Y_GE25","LT",2007,3.9,"Lithuania"
"Y_GE25","LT0",2007,3.9,"Lietuva"
"Y_GE25","LT00",2007,3.9,"Lietuva"
"Y_GE25","LU",2007,3.3,"Luxembourg"
"Y_GE25","LU0",2007,3.3,"Luxembourg"
"Y_GE25","LU00",2007,3.3,"Luxembourg"
"Y_GE25","LV",2007,5.4,"Latvia"
"Y_GE25","LV0",2007,5.4,"Latvija"
"Y_GE25","LV00",2007,5.4,"Latvija"
"Y_GE25","MK",2007,31.6,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2007,31.6,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2007,31.6,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2007,4.9,"Malta"
"Y_GE25","MT0",2007,4.9,"Malta"
"Y_GE25","MT00",2007,4.9,"Malta"
"Y_GE25","NL",2007,2.6,"Netherlands"
"Y_GE25","NL1",2007,3.1,"Noord-Nederland"
"Y_GE25","NL11",2007,3.9,"Groningen"
"Y_GE25","NL12",2007,2.6,"Friesland (NL)"
"Y_GE25","NL13",2007,3,"Drenthe"
"Y_GE25","NL2",2007,2.6,"Oost-Nederland"
"Y_GE25","NL21",2007,2.8,"Overijssel"
"Y_GE25","NL22",2007,2.3,"Gelderland"
"Y_GE25","NL23",2007,3.4,"Flevoland"
"Y_GE25","NL3",2007,2.6,"West-Nederland"
"Y_GE25","NL31",2007,2.2,"Utrecht"
"Y_GE25","NL32",2007,2.5,"Noord-Holland"
"Y_GE25","NL33",2007,2.9,"Zuid-Holland"
"Y_GE25","NL34",2007,1.5,"Zeeland"
"Y_GE25","NL4",2007,2.6,"Zuid-Nederland"
"Y_GE25","NL41",2007,2.3,"Noord-Brabant"
"Y_GE25","NL42",2007,3.3,"Limburg (NL)"
"Y_GE25","NO",2007,1.7,"Norway"
"Y_GE25","NO0",2007,1.7,"Norge"
"Y_GE25","NO01",2007,1.8,"Oslo og Akershus"
"Y_GE25","NO02",2007,1.2,"Hedmark og Oppland"
"Y_GE25","NO03",2007,2.1,"Sør-Østlandet"
"Y_GE25","NO04",2007,1.3,"Agder og Rogaland"
"Y_GE25","NO05",2007,1.5,"Vestlandet"
"Y_GE25","NO06",2007,2.1,"Trøndelag"
"Y_GE25","NO07",2007,1.7,"Nord-Norge"
"Y_GE25","PL",2007,8.1,"Poland"
"Y_GE25","PL1",2007,7.8,"Region Centralny"
"Y_GE25","PL11",2007,8.3,"Lódzkie"
"Y_GE25","PL12",2007,7.5,"Mazowieckie"
"Y_GE25","PL2",2007,6.8,"Region Poludniowy"
"Y_GE25","PL21",2007,6.4,"Malopolskie"
"Y_GE25","PL22",2007,7,"Slaskie"
"Y_GE25","PL3",2007,8.2,"Region Wschodni"
"Y_GE25","PL31",2007,7.6,"Lubelskie"
"Y_GE25","PL32",2007,7.8,"Podkarpackie"
"Y_GE25","PL33",2007,10.1,"Swietokrzyskie"
"Y_GE25","PL34",2007,7.6,"Podlaskie"
"Y_GE25","PL4",2007,7.9,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2007,6.7,"Wielkopolskie"
"Y_GE25","PL42",2007,10.2,"Zachodniopomorskie"
"Y_GE25","PL43",2007,8.3,"Lubuskie"
"Y_GE25","PL5",2007,10.6,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2007,11.4,"Dolnoslaskie"
"Y_GE25","PL52",2007,8.2,"Opolskie"
"Y_GE25","PL6",2007,8.9,"Region Pólnocny"
"Y_GE25","PL61",2007,9.7,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2007,9,"Warminsko-Mazurskie"
"Y_GE25","PL63",2007,7.9,"Pomorskie"
"Y_GE25","PT",2007,7.1,"Portugal"
"Y_GE25","PT1",2007,7.2,"Continente"
"Y_GE25","PT11",2007,8.5,"Norte"
"Y_GE25","PT15",2007,5.5,"Algarve"
"Y_GE25","PT16",2007,4.8,"Centro (PT)"
"Y_GE25","PT17",2007,8.1,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2007,7.2,"Alentejo"
"Y_GE25","PT2",2007,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2007,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2007,5.5,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2007,5.5,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2007,4.9,"Romania"
"Y_GE25","RO1",2007,4.9,"Macroregiunea unu"
"Y_GE25","RO11",2007,3.2,"Nord-Vest"
"Y_GE25","RO12",2007,6.7,"Centru"
"Y_GE25","RO2",2007,4.9,"Macroregiunea doi"
"Y_GE25","RO21",2007,3.9,"Nord-Est"
"Y_GE25","RO22",2007,6.4,"Sud-Est"
"Y_GE25","RO3",2007,5,"Macroregiunea trei"
"Y_GE25","RO31",2007,6.3,"Sud - Muntenia"
"Y_GE25","RO32",2007,3.1,"Bucuresti - Ilfov"
"Y_GE25","RO4",2007,4.9,"Macroregiunea patru"
"Y_GE25","RO41",2007,5.4,"Sud-Vest Oltenia"
"Y_GE25","RO42",2007,4.3,"Vest"
"Y_GE25","SE",2007,4.3,"Sweden"
"Y_GE25","SE1",2007,4.3,"Östra Sverige"
"Y_GE25","SE11",2007,3.9,"Stockholm"
"Y_GE25","SE12",2007,4.8,"Östra Mellansverige"
"Y_GE25","SE2",2007,4.1,"Södra Sverige"
"Y_GE25","SE21",2007,3.4,"Småland med öarna"
"Y_GE25","SE22",2007,4.8,"Sydsverige"
"Y_GE25","SE23",2007,3.9,"Västsverige"
"Y_GE25","SE3",2007,4.5,"Norra Sverige"
"Y_GE25","SE31",2007,4.4,"Norra Mellansverige"
"Y_GE25","SE32",2007,4.3,"Mellersta Norrland"
"Y_GE25","SE33",2007,4.9,"Övre Norrland"
"Y_GE25","SI",2007,4.2,"Slovenia"
"Y_GE25","SI0",2007,4.2,"Slovenija"
"Y_GE25","SI01",2007,4.8,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2007,3.5,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2007,10,"Slovakia"
"Y_GE25","SK0",2007,10,"Slovensko"
"Y_GE25","SK01",2007,4,"Bratislavský kraj"
"Y_GE25","SK02",2007,7.2,"Západné Slovensko"
"Y_GE25","SK03",2007,14.1,"Stredné Slovensko"
"Y_GE25","SK04",2007,12.9,"Východné Slovensko"
"Y_GE25","TR",2007,7,"Turkey"
"Y_GE25","TR1",2007,7.9,"Istanbul"
"Y_GE25","TR10",2007,7.9,"Istanbul"
"Y_GE25","TR2",2007,4.1,"Bati Marmara"
"Y_GE25","TR21",2007,4.7,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2007,3.5,"Balikesir, Çanakkale"
"Y_GE25","TR3",2007,6.4,"Ege"
"Y_GE25","TR31",2007,7.5,"Izmir"
"Y_GE25","TR32",2007,6.8,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2007,4.6,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2007,6.5,"Dogu Marmara"
"Y_GE25","TR41",2007,5.6,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2007,7.7,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2007,7.3,"Bati Anadolu"
"Y_GE25","TR51",2007,7.6,"Ankara"
"Y_GE25","TR52",2007,6.8,"Konya, Karaman"
"Y_GE25","TR6",2007,8,"Akdeniz"
"Y_GE25","TR61",2007,5.1,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2007,10.5,"Adana, Mersin"
"Y_GE25","TR63",2007,8,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2007,6,"Orta Anadolu"
"Y_GE25","TR71",2007,4.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2007,6.9,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2007,4.9,"Bati Karadeniz"
"Y_GE25","TR81",2007,4.5,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2007,2.2,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2007,5.7,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2007,3.1,"Dogu Karadeniz"
"Y_GE25","TR90",2007,3.1,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2007,3.6,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2007,3.5,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2007,3.7,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2007,8.3,"Ortadogu Anadolu"
"Y_GE25","TRB1",2007,7.6,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2007,9.2,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2007,13.5,"Güneydogu Anadolu"
"Y_GE25","TRC1",2007,15.1,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2007,10.7,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2007,15.4,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2007,3.6,"United Kingdom"
"Y_GE25","UKC",2007,4.1,"North East (UK)"
"Y_GE25","UKC1",2007,3.8,"Tees Valley and Durham"
"Y_GE25","UKC2",2007,4.4,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2007,4,"North West (UK)"
"Y_GE25","UKD1",2007,2.2,"Cumbria"
"Y_GE25","UKD3",2007,4.4,"Greater Manchester"
"Y_GE25","UKD4",2007,4,"Lancashire"
"Y_GE25","UKD6",2007,1.9,"Cheshire"
"Y_GE25","UKD7",2007,5.1,"Merseyside"
"Y_GE25","UKE",2007,3.8,"Yorkshire and The Humber"
"Y_GE25","UKE1",2007,4.2,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2007,2.4,"North Yorkshire"
"Y_GE25","UKE3",2007,4.6,"South Yorkshire"
"Y_GE25","UKE4",2007,3.6,"West Yorkshire"
"Y_GE25","UKF",2007,3.4,"East Midlands (UK)"
"Y_GE25","UKF1",2007,3.8,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2007,2.9,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2007,3.7,"Lincolnshire"
"Y_GE25","UKG",2007,4.4,"West Midlands (UK)"
"Y_GE25","UKG1",2007,2.9,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2007,3.6,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2007,5.7,"West Midlands"
"Y_GE25","UKH",2007,3.3,"East of England"
"Y_GE25","UKH1",2007,3,"East Anglia"
"Y_GE25","UKH2",2007,3.3,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2007,3.7,"Essex"
"Y_GE25","UKI",2007,4.9,"London"
"Y_GE25","UKI1",2007,6.2,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2007,4.1,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2007,3,"South East (UK)"
"Y_GE25","UKJ1",2007,2.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2007,2.6,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2007,3,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2007,3.7,"Kent"
"Y_GE25","UKK",2007,2.6,"South West (UK)"
"Y_GE25","UKK1",2007,2.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2007,2.4,"Dorset and Somerset"
"Y_GE25","UKK3",2007,3.4,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2007,2.8,"Devon"
"Y_GE25","UKL",2007,3.4,"Wales"
"Y_GE25","UKL1",2007,3.6,"West Wales and The Valleys"
"Y_GE25","UKL2",2007,3.2,"East Wales"
"Y_GE25","UKM",2007,3.2,"Scotland"
"Y_GE25","UKM2",2007,3.2,"Eastern Scotland"
"Y_GE25","UKM3",2007,3.6,"South Western Scotland"
"Y_GE25","UKM5",2007,2.4,"North Eastern Scotland"
"Y_GE25","UKM6",2007,NA,"Highlands and Islands"
"Y_GE25","UKN",2007,2.8,"Northern Ireland (UK)"
"Y_GE25","UKN0",2007,2.8,"Northern Ireland (UK)"
"Y15-24","AT",2006,9.8,"Austria"
"Y15-24","AT1",2006,13.7,"Ostösterreich"
"Y15-24","AT11",2006,NA,"Burgenland (AT)"
"Y15-24","AT12",2006,8.6,"Niederösterreich"
"Y15-24","AT13",2006,19.4,"Wien"
"Y15-24","AT2",2006,8.3,"Südösterreich"
"Y15-24","AT21",2006,8.6,"Kärnten"
"Y15-24","AT22",2006,8.2,"Steiermark"
"Y15-24","AT3",2006,6.8,"Westösterreich"
"Y15-24","AT31",2006,6.1,"Oberösterreich"
"Y15-24","AT32",2006,NA,"Salzburg"
"Y15-24","AT33",2006,6.7,"Tirol"
"Y15-24","AT34",2006,NA,"Vorarlberg"
"Y15-24","BE",2006,20.5,"Belgium"
"Y15-24","BE1",2006,35.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2006,35.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2006,12.5,"Vlaams Gewest"
"Y15-24","BE21",2006,13.4,"Prov. Antwerpen"
"Y15-24","BE22",2006,13.1,"Prov. Limburg (BE)"
"Y15-24","BE23",2006,10.9,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2006,14.8,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2006,10.9,"Prov. West-Vlaanderen"
"Y15-24","BE3",2006,31.3,"Région wallonne"
"Y15-24","BE31",2006,24.8,"Prov. Brabant Wallon"
"Y15-24","BE32",2006,36.8,"Prov. Hainaut"
"Y15-24","BE33",2006,30.6,"Prov. Liège"
"Y15-24","BE34",2006,23.8,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2006,28,"Prov. Namur"
"Y15-24","BG",2006,19.5,"Bulgaria"
"Y15-24","BG3",2006,23.3,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2006,25.8,"Severozapaden"
"Y15-24","BG32",2006,25.2,"Severen tsentralen"
"Y15-24","BG33",2006,23.6,"Severoiztochen"
"Y15-24","BG34",2006,19.3,"Yugoiztochen"
"Y15-24","BG4",2006,15.8,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2006,13,"Yugozapaden"
"Y15-24","BG42",2006,21.1,"Yuzhen tsentralen"
"Y15-24","CH",2006,7.7,"Switzerland"
"Y15-24","CH0",2006,7.7,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2006,10,"Région lémanique"
"Y15-24","CH02",2006,6.7,"Espace Mittelland"
"Y15-24","CH03",2006,8.6,"Nordwestschweiz"
"Y15-24","CH04",2006,8.1,"Zürich"
"Y15-24","CH05",2006,7.4,"Ostschweiz"
"Y15-24","CH06",2006,3.7,"Zentralschweiz"
"Y15-24","CH07",2006,12.1,"Ticino"
"Y15-24","CY",2006,10,"Cyprus"
"Y15-24","CY0",2006,10,"Kypros"
"Y15-24","CY00",2006,10,"Kypros"
"Y15-24","CZ",2006,17.5,"Czech Republic"
"Y15-24","CZ0",2006,17.5,"Ceská republika"
"Y15-24","CZ01",2006,8,"Praha"
"Y15-24","CZ02",2006,10.9,"Strední Cechy"
"Y15-24","CZ03",2006,11.4,"Jihozápad"
"Y15-24","CZ04",2006,28.1,"Severozápad"
"Y15-24","CZ05",2006,12,"Severovýchod"
"Y15-24","CZ06",2006,18.7,"Jihovýchod"
"Y15-24","CZ07",2006,15.3,"Strední Morava"
"Y15-24","CZ08",2006,30.5,"Moravskoslezsko"
"Y15-24","DE",2006,13.8,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2006,8.8,"Baden-Württemberg"
"Y15-24","DE11",2006,9.4,"Stuttgart"
"Y15-24","DE12",2006,9.7,"Karlsruhe"
"Y15-24","DE13",2006,6.4,"Freiburg"
"Y15-24","DE14",2006,9.5,"Tübingen"
"Y15-24","DE2",2006,8.6,"Bayern"
"Y15-24","DE21",2006,6.9,"Oberbayern"
"Y15-24","DE22",2006,11.1,"Niederbayern"
"Y15-24","DE23",2006,7.2,"Oberpfalz"
"Y15-24","DE24",2006,12,"Oberfranken"
"Y15-24","DE25",2006,8.8,"Mittelfranken"
"Y15-24","DE26",2006,10.2,"Unterfranken"
"Y15-24","DE27",2006,7.7,"Schwaben"
"Y15-24","DE3",2006,25.1,"Berlin"
"Y15-24","DE30",2006,25.1,"Berlin"
"Y15-24","DE4",2006,19.8,"Brandenburg"
"Y15-24","DE40",2006,19.8,"Brandenburg"
"Y15-24","DE5",2006,16.5,"Bremen"
"Y15-24","DE50",2006,16.5,"Bremen"
"Y15-24","DE6",2006,15.8,"Hamburg"
"Y15-24","DE60",2006,15.8,"Hamburg"
"Y15-24","DE7",2006,13.1,"Hessen"
"Y15-24","DE71",2006,12.5,"Darmstadt"
"Y15-24","DE72",2006,15.2,"Gießen"
"Y15-24","DE73",2006,12.5,"Kassel"
"Y15-24","DE8",2006,20.3,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2006,20.3,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2006,14.2,"Niedersachsen"
"Y15-24","DE91",2006,15,"Braunschweig"
"Y15-24","DE92",2006,13.5,"Hannover"
"Y15-24","DE93",2006,16.2,"Lüneburg"
"Y15-24","DE94",2006,13,"Weser-Ems"
"Y15-24","DEA",2006,14.4,"Nordrhein-Westfalen"
"Y15-24","DEA1",2006,14.5,"Düsseldorf"
"Y15-24","DEA2",2006,13.2,"Köln"
"Y15-24","DEA3",2006,15.1,"Münster"
"Y15-24","DEA4",2006,14.3,"Detmold"
"Y15-24","DEA5",2006,15,"Arnsberg"
"Y15-24","DEB",2006,13.3,"Rheinland-Pfalz"
"Y15-24","DEB1",2006,12.4,"Koblenz"
"Y15-24","DEB2",2006,NA,"Trier"
"Y15-24","DEB3",2006,15.4,"Rheinhessen-Pfalz"
"Y15-24","DEC",2006,13.9,"Saarland"
"Y15-24","DEC0",2006,13.9,"Saarland"
"Y15-24","DED",2006,18.4,"Sachsen"
"Y15-24","DED2",2006,19.5,"Dresden"
"Y15-24","DED4",2006,16.8,"Chemnitz"
"Y15-24","DED5",2006,18.8,"Leipzig"
"Y15-24","DEE",2006,18.9,"Sachsen-Anhalt"
"Y15-24","DEE0",2006,18.9,"Sachsen-Anhalt"
"Y15-24","DEF",2006,13.3,"Schleswig-Holstein"
"Y15-24","DEF0",2006,13.3,"Schleswig-Holstein"
"Y15-24","DEG",2006,17.4,"Thüringen"
"Y15-24","DEG0",2006,17.4,"Thüringen"
"Y15-24","DK",2006,7.7,"Denmark"
"Y15-24","DK0",2006,7.7,"Danmark"
"Y15-24","EA17",2006,16.8,"Euro area (17 countries)"
"Y15-24","EA18",2006,16.8,"Euro area (18 countries)"
"Y15-24","EA19",2006,16.7,"Euro area (19 countries)"
"Y15-24","EE",2006,12.1,"Estonia"
"Y15-24","EE0",2006,12.1,"Eesti"
"Y15-24","EE00",2006,12.1,"Eesti"
"Y15-24","EL",2006,25,"Greece"
"Y15-24","EL1",2006,27,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2006,31.3,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2006,26.6,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2006,28,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2006,23.9,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2006,30.2,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2006,32.5,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2006,32.3,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2006,33.6,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2006,26.8,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2006,27.3,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2006,21.5,"Attiki"
"Y15-24","EL30",2006,21.5,"Attiki"
"Y15-24","EL4",2006,21.2,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2006,34.9,"Voreio Aigaio"
"Y15-24","EL42",2006,17.9,"Notio Aigaio"
"Y15-24","EL43",2006,18.7,"Kriti"
"Y15-24","ES",2006,17.9,"Spain"
"Y15-24","ES1",2006,18.7,"Noroeste (ES)"
"Y15-24","ES11",2006,17.8,"Galicia"
"Y15-24","ES12",2006,22.4,"Principado de Asturias"
"Y15-24","ES13",2006,16.7,"Cantabria"
"Y15-24","ES2",2006,16.6,"Noreste (ES)"
"Y15-24","ES21",2006,21.1,"País Vasco"
"Y15-24","ES22",2006,14.2,"Comunidad Foral de Navarra"
"Y15-24","ES23",2006,14.9,"La Rioja"
"Y15-24","ES24",2006,11.8,"Aragón"
"Y15-24","ES3",2006,14.7,"Comunidad de Madrid"
"Y15-24","ES30",2006,14.7,"Comunidad de Madrid"
"Y15-24","ES4",2006,18.4,"Centro (ES)"
"Y15-24","ES41",2006,16.9,"Castilla y León"
"Y15-24","ES42",2006,17,"Castilla-la Mancha"
"Y15-24","ES43",2006,24.2,"Extremadura"
"Y15-24","ES5",2006,15.8,"Este (ES)"
"Y15-24","ES51",2006,14.6,"Cataluña"
"Y15-24","ES52",2006,17.9,"Comunidad Valenciana"
"Y15-24","ES53",2006,13.4,"Illes Balears"
"Y15-24","ES6",2006,21.2,"Sur (ES)"
"Y15-24","ES61",2006,21.7,"Andalucía"
"Y15-24","ES62",2006,17.1,"Región de Murcia"
"Y15-24","ES63",2006,54.8,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2006,23.7,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2006,23.4,"Canarias (ES)"
"Y15-24","ES70",2006,23.4,"Canarias (ES)"
"Y15-24","EU15",2006,16.1,"European Union (15 countries)"
"Y15-24","EU27",2006,17.4,"European Union (27 countries)"
"Y15-24","EU28",2006,17.5,"European Union (28 countries)"
"Y15-24","FI",2006,18.7,"Finland"
"Y15-24","FI1",2006,18.7,"Manner-Suomi"
"Y15-24","FI19",2006,19,"Länsi-Suomi"
"Y15-24","FI1B",2006,14.2,"Helsinki-Uusimaa"
"Y15-24","FI1C",2006,17.1,"Etelä-Suomi"
"Y15-24","FI1D",2006,25.7,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2006,NA,"Åland"
"Y15-24","FI20",2006,NA,"Åland"
"Y15-24","FR",2006,22.3,"France"
"Y15-24","FR1",2006,20,"Île de France"
"Y15-24","FR10",2006,20,"Île de France"
"Y15-24","FR2",2006,22.6,"Bassin Parisien"
"Y15-24","FR21",2006,18.3,"Champagne-Ardenne"
"Y15-24","FR22",2006,27.9,"Picardie"
"Y15-24","FR23",2006,25.5,"Haute-Normandie"
"Y15-24","FR24",2006,20.3,"Centre (FR)"
"Y15-24","FR25",2006,22.6,"Basse-Normandie"
"Y15-24","FR26",2006,19.3,"Bourgogne"
"Y15-24","FR3",2006,28.1,"Nord - Pas-de-Calais"
"Y15-24","FR30",2006,28.1,"Nord - Pas-de-Calais"
"Y15-24","FR4",2006,21.1,"Est (FR)"
"Y15-24","FR41",2006,24.6,"Lorraine"
"Y15-24","FR42",2006,16,"Alsace"
"Y15-24","FR43",2006,20.6,"Franche-Comté"
"Y15-24","FR5",2006,18.6,"Ouest (FR)"
"Y15-24","FR51",2006,17.5,"Pays de la Loire"
"Y15-24","FR52",2006,18.7,"Bretagne"
"Y15-24","FR53",2006,20.7,"Poitou-Charentes"
"Y15-24","FR6",2006,17.3,"Sud-Ouest (FR)"
"Y15-24","FR61",2006,19.4,"Aquitaine"
"Y15-24","FR62",2006,14.6,"Midi-Pyrénées"
"Y15-24","FR63",2006,NA,"Limousin"
"Y15-24","FR7",2006,19.2,"Centre-Est (FR)"
"Y15-24","FR71",2006,19.5,"Rhône-Alpes"
"Y15-24","FR72",2006,18,"Auvergne"
"Y15-24","FR8",2006,26.7,"Méditerranée"
"Y15-24","FR81",2006,27.9,"Languedoc-Roussillon"
"Y15-24","FR82",2006,26.1,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2006,NA,"Corse"
"Y15-24","FR9",2006,52.9,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2006,59.9,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2006,56.1,"Martinique (NUTS 2010)"
"Y15-24","FR93",2006,49.4,"Guyane (NUTS 2010)"
"Y15-24","FR94",2006,50.4,"Réunion (NUTS 2010)"
"Y15-24","HR",2006,28.9,"Croatia"
"Y15-24","HR0",2006,28.9,"Hrvatska"
"Y15-24","HU",2006,19.1,"Hungary"
"Y15-24","HU1",2006,14.8,"Közép-Magyarország"
"Y15-24","HU10",2006,14.8,"Közép-Magyarország"
"Y15-24","HU2",2006,15.9,"Dunántúl"
"Y15-24","HU21",2006,13.3,"Közép-Dunántúl"
"Y15-24","HU22",2006,13.5,"Nyugat-Dunántúl"
"Y15-24","HU23",2006,22.5,"Dél-Dunántúl"
"Y15-24","HU3",2006,24.5,"Alföld és Észak"
"Y15-24","HU31",2006,25.9,"Észak-Magyarország"
"Y15-24","HU32",2006,26.6,"Észak-Alföld"
"Y15-24","HU33",2006,20.4,"Dél-Alföld"
"Y15-24","IE",2006,8.6,"Ireland"
"Y15-24","IE0",2006,8.6,"Éire/Ireland"
"Y15-24","IE01",2006,9.9,"Border, Midland and Western"
"Y15-24","IE02",2006,8.1,"Southern and Eastern"
"Y15-24","IS",2006,8.3,"Iceland"
"Y15-24","IS0",2006,8.3,"Ísland"
"Y15-24","IS00",2006,8.3,"Ísland"
"Y15-24","IT",2006,21.8,"Italy"
"Y15-24","ITC",2006,13.6,"Nord-Ovest"
"Y15-24","ITC1",2006,15.7,"Piemonte"
"Y15-24","ITC2",2006,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2006,16.4,"Liguria"
"Y15-24","ITC4",2006,12.4,"Lombardia"
"Y15-24","ITF",2006,33.1,"Sud"
"Y15-24","ITF1",2006,21.1,"Abruzzo"
"Y15-24","ITF2",2006,28,"Molise"
"Y15-24","ITF3",2006,35.8,"Campania"
"Y15-24","ITF4",2006,32.3,"Puglia"
"Y15-24","ITF5",2006,31.9,"Basilicata"
"Y15-24","ITF6",2006,35.1,"Calabria"
"Y15-24","ITG",2006,36.9,"Isole"
"Y15-24","ITG1",2006,38.9,"Sicilia"
"Y15-24","ITG2",2006,31.1,"Sardegna"
"Y15-24","ITH",2006,11,"Nord-Est"
"Y15-24","ITH1",2006,7.2,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2006,9.4,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2006,11.8,"Veneto"
"Y15-24","ITH4",2006,11.5,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2006,10.7,"Emilia-Romagna"
"Y15-24","ITI",2006,19.8,"Centro (IT)"
"Y15-24","ITI1",2006,15.8,"Toscana"
"Y15-24","ITI2",2006,14.6,"Umbria"
"Y15-24","ITI3",2006,11.9,"Marche"
"Y15-24","ITI4",2006,26.1,"Lazio"
"Y15-24","LT",2006,10,"Lithuania"
"Y15-24","LT0",2006,10,"Lietuva"
"Y15-24","LT00",2006,10,"Lietuva"
"Y15-24","LU",2006,16.2,"Luxembourg"
"Y15-24","LU0",2006,16.2,"Luxembourg"
"Y15-24","LU00",2006,16.2,"Luxembourg"
"Y15-24","LV",2006,13.6,"Latvia"
"Y15-24","LV0",2006,13.6,"Latvija"
"Y15-24","LV00",2006,13.6,"Latvija"
"Y15-24","MK",2006,59.7,"Former Yugoslav Republic of Macedonia, the"
"Y15-24","MK0",2006,59.7,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MK00",2006,59.7,"Poranesna jugoslovenska Republika Makedonija"
"Y15-24","MT",2006,15.5,"Malta"
"Y15-24","MT0",2006,15.5,"Malta"
"Y15-24","MT00",2006,15.5,"Malta"
"Y15-24","NL",2006,6.6,"Netherlands"
"Y15-24","NL1",2006,8,"Noord-Nederland"
"Y15-24","NL11",2006,8.1,"Groningen"
"Y15-24","NL12",2006,7.1,"Friesland (NL)"
"Y15-24","NL13",2006,9.4,"Drenthe"
"Y15-24","NL2",2006,6,"Oost-Nederland"
"Y15-24","NL21",2006,6,"Overijssel"
"Y15-24","NL22",2006,5.2,"Gelderland"
"Y15-24","NL23",2006,10,"Flevoland"
"Y15-24","NL3",2006,6.8,"West-Nederland"
"Y15-24","NL31",2006,5.8,"Utrecht"
"Y15-24","NL32",2006,6.5,"Noord-Holland"
"Y15-24","NL33",2006,7.7,"Zuid-Holland"
"Y15-24","NL34",2006,NA,"Zeeland"
"Y15-24","NL4",2006,5.9,"Zuid-Nederland"
"Y15-24","NL41",2006,5,"Noord-Brabant"
"Y15-24","NL42",2006,8,"Limburg (NL)"
"Y15-24","NO",2006,8.7,"Norway"
"Y15-24","NO0",2006,8.7,"Norge"
"Y15-24","NO01",2006,7.8,"Oslo og Akershus"
"Y15-24","NO02",2006,10,"Hedmark og Oppland"
"Y15-24","NO03",2006,10.7,"Sør-Østlandet"
"Y15-24","NO04",2006,6.8,"Agder og Rogaland"
"Y15-24","NO05",2006,7.7,"Vestlandet"
"Y15-24","NO06",2006,10,"Trøndelag"
"Y15-24","NO07",2006,10.1,"Nord-Norge"
"Y15-24","PL",2006,29.8,"Poland"
"Y15-24","PL1",2006,27.3,"Region Centralny"
"Y15-24","PL11",2006,25,"Lódzkie"
"Y15-24","PL12",2006,28.6,"Mazowieckie"
"Y15-24","PL2",2006,30,"Region Poludniowy"
"Y15-24","PL21",2006,30.2,"Malopolskie"
"Y15-24","PL22",2006,29.8,"Slaskie"
"Y15-24","PL3",2006,33.7,"Region Wschodni"
"Y15-24","PL31",2006,32.1,"Lubelskie"
"Y15-24","PL32",2006,35.3,"Podkarpackie"
"Y15-24","PL33",2006,36.6,"Swietokrzyskie"
"Y15-24","PL34",2006,29.9,"Podlaskie"
"Y15-24","PL4",2006,28.6,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2006,27.1,"Wielkopolskie"
"Y15-24","PL42",2006,32.4,"Zachodniopomorskie"
"Y15-24","PL43",2006,29.3,"Lubuskie"
"Y15-24","PL5",2006,31.9,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2006,32.8,"Dolnoslaskie"
"Y15-24","PL52",2006,29.1,"Opolskie"
"Y15-24","PL6",2006,30.2,"Region Pólnocny"
"Y15-24","PL61",2006,31.1,"Kujawsko-Pomorskie"
"Y15-24","PL62",2006,33.5,"Warminsko-Mazurskie"
"Y15-24","PL63",2006,27.3,"Pomorskie"
"Y15-24","PT",2006,16.5,"Portugal"
"Y15-24","PT1",2006,16.9,"Continente"
"Y15-24","PT11",2006,17,"Norte"
"Y15-24","PT15",2006,NA,"Algarve"
"Y15-24","PT16",2006,12.2,"Centro (PT)"
"Y15-24","PT17",2006,19.8,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2006,21.1,"Alentejo"
"Y15-24","PT2",2006,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2006,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2006,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2006,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2006,21.4,"Romania"
"Y15-24","RO1",2006,20.6,"Macroregiunea unu"
"Y15-24","RO11",2006,18.6,"Nord-Vest"
"Y15-24","RO12",2006,22.7,"Centru"
"Y15-24","RO2",2006,21,"Macroregiunea doi"
"Y15-24","RO21",2006,18.1,"Nord-Est"
"Y15-24","RO22",2006,24.8,"Sud-Est"
"Y15-24","RO3",2006,23.7,"Macroregiunea trei"
"Y15-24","RO31",2006,27,"Sud - Muntenia"
"Y15-24","RO32",2006,15.9,"Bucuresti - Ilfov"
"Y15-24","RO4",2006,19.9,"Macroregiunea patru"
"Y15-24","RO41",2006,23.4,"Sud-Vest Oltenia"
"Y15-24","RO42",2006,15.8,"Vest"
"Y15-24","SE",2006,21.5,"Sweden"
"Y15-24","SE1",2006,21.1,"Östra Sverige"
"Y15-24","SE11",2006,19.5,"Stockholm"
"Y15-24","SE12",2006,23.1,"Östra Mellansverige"
"Y15-24","SE2",2006,21.3,"Södra Sverige"
"Y15-24","SE21",2006,17.6,"Småland med öarna"
"Y15-24","SE22",2006,25.1,"Sydsverige"
"Y15-24","SE23",2006,20.4,"Västsverige"
"Y15-24","SE3",2006,22.7,"Norra Sverige"
"Y15-24","SE31",2006,23.8,"Norra Mellansverige"
"Y15-24","SE32",2006,19.4,"Mellersta Norrland"
"Y15-24","SE33",2006,23.1,"Övre Norrland"
"Y15-24","SI",2006,13.9,"Slovenia"
"Y15-24","SI0",2006,13.9,"Slovenija"
"Y15-24","SI01",2006,17.1,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2006,10.1,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2006,26.6,"Slovakia"
"Y15-24","SK0",2006,26.6,"Slovensko"
"Y15-24","SK01",2006,8,"Bratislavský kraj"
"Y15-24","SK02",2006,21.9,"Západné Slovensko"
"Y15-24","SK03",2006,28.8,"Stredné Slovensko"
"Y15-24","SK04",2006,35.7,"Východné Slovensko"
"Y15-24","TR",2006,16.4,"Turkey"
"Y15-24","TR1",2006,16.1,"Istanbul"
"Y15-24","TR10",2006,16.1,"Istanbul"
"Y15-24","TR2",2006,14.5,"Bati Marmara"
"Y15-24","TR21",2006,15.3,"Tekirdag, Edirne, Kirklareli"
"Y15-24","TR22",2006,13.4,"Balikesir, Çanakkale"
"Y15-24","TR3",2006,14.3,"Ege"
"Y15-24","TR31",2006,17.8,"Izmir"
"Y15-24","TR32",2006,10.7,"Aydin, Denizli, Mugla"
"Y15-24","TR33",2006,13,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y15-24","TR4",2006,16.7,"Dogu Marmara"
"Y15-24","TR41",2006,15,"Bursa, Eskisehir, Bilecik"
"Y15-24","TR42",2006,18.8,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y15-24","TR5",2006,22,"Bati Anadolu"
"Y15-24","TR51",2006,23.3,"Ankara"
"Y15-24","TR52",2006,19.2,"Konya, Karaman"
"Y15-24","TR6",2006,17.6,"Akdeniz"
"Y15-24","TR61",2006,11.8,"Antalya, Isparta, Burdur"
"Y15-24","TR62",2006,24.8,"Adana, Mersin"
"Y15-24","TR63",2006,13.9,"Hatay, Kahramanmaras, Osmaniye"
"Y15-24","TR7",2006,21.5,"Orta Anadolu"
"Y15-24","TR71",2006,19.1,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y15-24","TR72",2006,23.7,"Kayseri, Sivas, Yozgat"
"Y15-24","TR8",2006,11.5,"Bati Karadeniz"
"Y15-24","TR81",2006,13.4,"Zonguldak, Karabük, Bartin"
"Y15-24","TR82",2006,10.5,"Kastamonu, Çankiri, Sinop"
"Y15-24","TR83",2006,11,"Samsun, Tokat, Çorum, Amasya"
"Y15-24","TR9",2006,13.5,"Dogu Karadeniz"
"Y15-24","TR90",2006,13.5,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y15-24","TRA",2006,8.4,"Kuzeydogu Anadolu"
"Y15-24","TRA1",2006,7.7,"Erzurum, Erzincan, Bayburt"
"Y15-24","TRA2",2006,9.1,"Agri, Kars, Igdir, Ardahan"
"Y15-24","TRB",2006,17.9,"Ortadogu Anadolu"
"Y15-24","TRB1",2006,25.7,"Malatya, Elazig, Bingöl, Tunceli"
"Y15-24","TRB2",2006,11.4,"Van, Mus, Bitlis, Hakkari"
"Y15-24","TRC",2006,19,"Güneydogu Anadolu"
"Y15-24","TRC1",2006,17.4,"Gaziantep, Adiyaman, Kilis"
"Y15-24","TRC2",2006,17.9,"Sanliurfa, Diyarbakir"
"Y15-24","TRC3",2006,24.7,"Mardin, Batman, Sirnak, Siirt"
"Y15-24","UK",2006,13.9,"United Kingdom"
"Y15-24","UKC",2006,15,"North East (UK)"
"Y15-24","UKC1",2006,15.6,"Tees Valley and Durham"
"Y15-24","UKC2",2006,14.5,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2006,13.7,"North West (UK)"
"Y15-24","UKD1",2006,11.6,"Cumbria"
"Y15-24","UKD3",2006,12.8,"Greater Manchester"
"Y15-24","UKD4",2006,14.8,"Lancashire"
"Y15-24","UKD6",2006,9.1,"Cheshire"
"Y15-24","UKD7",2006,17.2,"Merseyside"
"Y15-24","UKE",2006,14.8,"Yorkshire and The Humber"
"Y15-24","UKE1",2006,14.7,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2006,13.1,"North Yorkshire"
"Y15-24","UKE3",2006,16.9,"South Yorkshire"
"Y15-24","UKE4",2006,14.2,"West Yorkshire"
"Y15-24","UKF",2006,14.7,"East Midlands (UK)"
"Y15-24","UKF1",2006,15.7,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2006,14.5,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2006,12.3,"Lincolnshire"
"Y15-24","UKG",2006,16,"West Midlands (UK)"
"Y15-24","UKG1",2006,12.5,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2006,13,"Shropshire and Staffordshire"
"Y15-24","UKG3",2006,18.9,"West Midlands"
"Y15-24","UKH",2006,12.2,"East of England"
"Y15-24","UKH1",2006,12.4,"East Anglia"
"Y15-24","UKH2",2006,13.1,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2006,11.2,"Essex"
"Y15-24","UKI",2006,19.5,"London"
"Y15-24","UKI1",2006,20.3,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2006,18.9,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2006,11.6,"South East (UK)"
"Y15-24","UKJ1",2006,11.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2006,9.8,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2006,11.1,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2006,15.1,"Kent"
"Y15-24","UKK",2006,9.9,"South West (UK)"
"Y15-24","UKK1",2006,9.2,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2006,7.5,"Dorset and Somerset"
"Y15-24","UKK3",2006,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2006,14.2,"Devon"
"Y15-24","UKL",2006,13.6,"Wales"
"Y15-24","UKL1",2006,15,"West Wales and The Valleys"
"Y15-24","UKL2",2006,11.4,"East Wales"
"Y15-24","UKM",2006,13.5,"Scotland"
"Y15-24","UKM2",2006,15.7,"Eastern Scotland"
"Y15-24","UKM3",2006,13.4,"South Western Scotland"
"Y15-24","UKM5",2006,NA,"North Eastern Scotland"
"Y15-24","UKM6",2006,NA,"Highlands and Islands"
"Y15-24","UKN",2006,9.8,"Northern Ireland (UK)"
"Y15-24","UKN0",2006,9.8,"Northern Ireland (UK)"
"Y20-64","AT",2006,4.9,"Austria"
"Y20-64","AT1",2006,6.6,"Ostösterreich"
"Y20-64","AT11",2006,5,"Burgenland (AT)"
"Y20-64","AT12",2006,4.1,"Niederösterreich"
"Y20-64","AT13",2006,9.1,"Wien"
"Y20-64","AT2",2006,4.2,"Südösterreich"
"Y20-64","AT21",2006,4.5,"Kärnten"
"Y20-64","AT22",2006,4.1,"Steiermark"
"Y20-64","AT3",2006,3.3,"Westösterreich"
"Y20-64","AT31",2006,3.3,"Oberösterreich"
"Y20-64","AT32",2006,3.2,"Salzburg"
"Y20-64","AT33",2006,2.8,"Tirol"
"Y20-64","AT34",2006,4.6,"Vorarlberg"
"Y20-64","BE",2006,8,"Belgium"
"Y20-64","BE1",2006,17.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2006,17.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2006,4.8,"Vlaams Gewest"
"Y20-64","BE21",2006,5.6,"Prov. Antwerpen"
"Y20-64","BE22",2006,5.9,"Prov. Limburg (BE)"
"Y20-64","BE23",2006,4.4,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2006,4,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2006,3.9,"Prov. West-Vlaanderen"
"Y20-64","BE3",2006,11.4,"Région wallonne"
"Y20-64","BE31",2006,7.4,"Prov. Brabant Wallon"
"Y20-64","BE32",2006,14.1,"Prov. Hainaut"
"Y20-64","BE33",2006,11.3,"Prov. Liège"
"Y20-64","BE34",2006,7.6,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2006,10.2,"Prov. Namur"
"Y20-64","BG",2006,8.6,"Bulgaria"
"Y20-64","BG3",2006,10.4,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2006,10.7,"Severozapaden"
"Y20-64","BG32",2006,12.9,"Severen tsentralen"
"Y20-64","BG33",2006,10.5,"Severoiztochen"
"Y20-64","BG34",2006,7.8,"Yugoiztochen"
"Y20-64","BG4",2006,6.9,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2006,6.2,"Yugozapaden"
"Y20-64","BG42",2006,7.9,"Yuzhen tsentralen"
"Y20-64","CH",2006,3.8,"Switzerland"
"Y20-64","CH0",2006,3.8,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2006,4.9,"Région lémanique"
"Y20-64","CH02",2006,3.6,"Espace Mittelland"
"Y20-64","CH03",2006,3.9,"Nordwestschweiz"
"Y20-64","CH04",2006,3.5,"Zürich"
"Y20-64","CH05",2006,3.7,"Ostschweiz"
"Y20-64","CH06",2006,2.6,"Zentralschweiz"
"Y20-64","CH07",2006,5.2,"Ticino"
"Y20-64","CY",2006,4.5,"Cyprus"
"Y20-64","CY0",2006,4.5,"Kypros"
"Y20-64","CY00",2006,4.5,"Kypros"
"Y20-64","CZ",2006,6.9,"Czech Republic"
"Y20-64","CZ0",2006,6.9,"Ceská republika"
"Y20-64","CZ01",2006,2.8,"Praha"
"Y20-64","CZ02",2006,4.4,"Strední Cechy"
"Y20-64","CZ03",2006,4.6,"Jihozápad"
"Y20-64","CZ04",2006,12,"Severozápad"
"Y20-64","CZ05",2006,5.8,"Severovýchod"
"Y20-64","CZ06",2006,6.9,"Jihovýchod"
"Y20-64","CZ07",2006,7.5,"Strední Morava"
"Y20-64","CZ08",2006,11.5,"Moravskoslezsko"
"Y20-64","DE",2006,10.2,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2006,6.3,"Baden-Württemberg"
"Y20-64","DE11",2006,6.4,"Stuttgart"
"Y20-64","DE12",2006,7.2,"Karlsruhe"
"Y20-64","DE13",2006,5.5,"Freiburg"
"Y20-64","DE14",2006,5.8,"Tübingen"
"Y20-64","DE2",2006,6.4,"Bayern"
"Y20-64","DE21",2006,5.3,"Oberbayern"
"Y20-64","DE22",2006,6.4,"Niederbayern"
"Y20-64","DE23",2006,6.9,"Oberpfalz"
"Y20-64","DE24",2006,9.3,"Oberfranken"
"Y20-64","DE25",2006,7.9,"Mittelfranken"
"Y20-64","DE26",2006,6,"Unterfranken"
"Y20-64","DE27",2006,6.1,"Schwaben"
"Y20-64","DE3",2006,18.6,"Berlin"
"Y20-64","DE30",2006,18.6,"Berlin"
"Y20-64","DE4",2006,16.7,"Brandenburg"
"Y20-64","DE40",2006,16.7,"Brandenburg"
"Y20-64","DE5",2006,14.5,"Bremen"
"Y20-64","DE50",2006,14.5,"Bremen"
"Y20-64","DE6",2006,9.7,"Hamburg"
"Y20-64","DE60",2006,9.7,"Hamburg"
"Y20-64","DE7",2006,8,"Hessen"
"Y20-64","DE71",2006,7.9,"Darmstadt"
"Y20-64","DE72",2006,8.2,"Gießen"
"Y20-64","DE73",2006,8.5,"Kassel"
"Y20-64","DE8",2006,19.6,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2006,19.6,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2006,9.7,"Niedersachsen"
"Y20-64","DE91",2006,10.1,"Braunschweig"
"Y20-64","DE92",2006,10.5,"Hannover"
"Y20-64","DE93",2006,8.8,"Lüneburg"
"Y20-64","DE94",2006,9.3,"Weser-Ems"
"Y20-64","DEA",2006,9.7,"Nordrhein-Westfalen"
"Y20-64","DEA1",2006,9.6,"Düsseldorf"
"Y20-64","DEA2",2006,9,"Köln"
"Y20-64","DEA3",2006,9,"Münster"
"Y20-64","DEA4",2006,9.9,"Detmold"
"Y20-64","DEA5",2006,11,"Arnsberg"
"Y20-64","DEB",2006,7.9,"Rheinland-Pfalz"
"Y20-64","DEB1",2006,7.5,"Koblenz"
"Y20-64","DEB2",2006,6.3,"Trier"
"Y20-64","DEB3",2006,8.5,"Rheinhessen-Pfalz"
"Y20-64","DEC",2006,9.3,"Saarland"
"Y20-64","DEC0",2006,9.3,"Saarland"
"Y20-64","DED",2006,16.9,"Sachsen"
"Y20-64","DED2",2006,16.4,"Dresden"
"Y20-64","DED4",2006,16.8,"Chemnitz"
"Y20-64","DED5",2006,17.7,"Leipzig"
"Y20-64","DEE",2006,18,"Sachsen-Anhalt"
"Y20-64","DEE0",2006,18,"Sachsen-Anhalt"
"Y20-64","DEF",2006,8.9,"Schleswig-Holstein"
"Y20-64","DEF0",2006,8.9,"Schleswig-Holstein"
"Y20-64","DEG",2006,15.9,"Thüringen"
"Y20-64","DEG0",2006,15.9,"Thüringen"
"Y20-64","DK",2006,3.5,"Denmark"
"Y20-64","DK0",2006,3.5,"Danmark"
"Y20-64","EA17",2006,8.1,"Euro area (17 countries)"
"Y20-64","EA18",2006,8.1,"Euro area (18 countries)"
"Y20-64","EA19",2006,8.1,"Euro area (19 countries)"
"Y20-64","EE",2006,5.7,"Estonia"
"Y20-64","EE0",2006,5.7,"Eesti"
"Y20-64","EE00",2006,5.7,"Eesti"
"Y20-64","EL",2006,8.9,"Greece"
"Y20-64","EL1",2006,9.7,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2006,10.7,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2006,9.2,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2006,14.4,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2006,8.4,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2006,9.1,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2006,9.7,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2006,11.2,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2006,9.4,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2006,9,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2006,7.6,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2006,8.3,"Attiki"
"Y20-64","EL30",2006,8.3,"Attiki"
"Y20-64","EL4",2006,8,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2006,9.2,"Voreio Aigaio"
"Y20-64","EL42",2006,8.9,"Notio Aigaio"
"Y20-64","EL43",2006,7.2,"Kriti"
"Y20-64","ES",2006,8,"Spain"
"Y20-64","ES1",2006,8.1,"Noroeste (ES)"
"Y20-64","ES11",2006,8.2,"Galicia"
"Y20-64","ES12",2006,9,"Principado de Asturias"
"Y20-64","ES13",2006,6.2,"Cantabria"
"Y20-64","ES2",2006,6,"Noreste (ES)"
"Y20-64","ES21",2006,6.7,"País Vasco"
"Y20-64","ES22",2006,5.2,"Comunidad Foral de Navarra"
"Y20-64","ES23",2006,5.8,"La Rioja"
"Y20-64","ES24",2006,5.2,"Aragón"
"Y20-64","ES3",2006,5.8,"Comunidad de Madrid"
"Y20-64","ES30",2006,5.8,"Comunidad de Madrid"
"Y20-64","ES4",2006,8.9,"Centro (ES)"
"Y20-64","ES41",2006,7.8,"Castilla y León"
"Y20-64","ES42",2006,8.3,"Castilla-la Mancha"
"Y20-64","ES43",2006,12.6,"Extremadura"
"Y20-64","ES5",2006,6.6,"Este (ES)"
"Y20-64","ES51",2006,6.1,"Cataluña"
"Y20-64","ES52",2006,7.7,"Comunidad Valenciana"
"Y20-64","ES53",2006,5.9,"Illes Balears"
"Y20-64","ES6",2006,11.4,"Sur (ES)"
"Y20-64","ES61",2006,12,"Andalucía"
"Y20-64","ES62",2006,7.3,"Región de Murcia"
"Y20-64","ES63",2006,19.6,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2006,12.8,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2006,10.9,"Canarias (ES)"
"Y20-64","ES70",2006,10.9,"Canarias (ES)"
"Y20-64","EU15",2006,7.4,"European Union (15 countries)"
"Y20-64","EU27",2006,7.9,"European Union (27 countries)"
"Y20-64","EU28",2006,7.9,"European Union (28 countries)"
"Y20-64","FI",2006,7,"Finland"
"Y20-64","FI1",2006,7,"Manner-Suomi"
"Y20-64","FI19",2006,7.1,"Länsi-Suomi"
"Y20-64","FI1B",2006,4.7,"Helsinki-Uusimaa"
"Y20-64","FI1C",2006,7.1,"Etelä-Suomi"
"Y20-64","FI1D",2006,9.9,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2006,NA,"Åland"
"Y20-64","FI20",2006,NA,"Åland"
"Y20-64","FR",2006,8.5,"France"
"Y20-64","FR1",2006,8.2,"Île de France"
"Y20-64","FR10",2006,8.2,"Île de France"
"Y20-64","FR2",2006,7.5,"Bassin Parisien"
"Y20-64","FR21",2006,6.5,"Champagne-Ardenne"
"Y20-64","FR22",2006,9.6,"Picardie"
"Y20-64","FR23",2006,8,"Haute-Normandie"
"Y20-64","FR24",2006,6.4,"Centre (FR)"
"Y20-64","FR25",2006,6.7,"Basse-Normandie"
"Y20-64","FR26",2006,8.2,"Bourgogne"
"Y20-64","FR3",2006,11.3,"Nord - Pas-de-Calais"
"Y20-64","FR30",2006,11.3,"Nord - Pas-de-Calais"
"Y20-64","FR4",2006,7.3,"Est (FR)"
"Y20-64","FR41",2006,8.6,"Lorraine"
"Y20-64","FR42",2006,6,"Alsace"
"Y20-64","FR43",2006,6.9,"Franche-Comté"
"Y20-64","FR5",2006,6.8,"Ouest (FR)"
"Y20-64","FR51",2006,6.5,"Pays de la Loire"
"Y20-64","FR52",2006,7,"Bretagne"
"Y20-64","FR53",2006,7.1,"Poitou-Charentes"
"Y20-64","FR6",2006,7.2,"Sud-Ouest (FR)"
"Y20-64","FR61",2006,7.1,"Aquitaine"
"Y20-64","FR62",2006,7.7,"Midi-Pyrénées"
"Y20-64","FR63",2006,5.6,"Limousin"
"Y20-64","FR7",2006,7,"Centre-Est (FR)"
"Y20-64","FR71",2006,6.9,"Rhône-Alpes"
"Y20-64","FR72",2006,7.1,"Auvergne"
"Y20-64","FR8",2006,10.5,"Méditerranée"
"Y20-64","FR81",2006,10.4,"Languedoc-Roussillon"
"Y20-64","FR82",2006,10.5,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2006,10.7,"Corse"
"Y20-64","FR9",2006,26.1,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2006,26.6,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2006,23.5,"Martinique (NUTS 2010)"
"Y20-64","FR93",2006,27.8,"Guyane (NUTS 2010)"
"Y20-64","FR94",2006,26.9,"Réunion (NUTS 2010)"
"Y20-64","HR",2006,10.8,"Croatia"
"Y20-64","HR0",2006,10.8,"Hrvatska"
"Y20-64","HU",2006,7.3,"Hungary"
"Y20-64","HU1",2006,5,"Közép-Magyarország"
"Y20-64","HU10",2006,5,"Közép-Magyarország"
"Y20-64","HU2",2006,6.7,"Dunántúl"
"Y20-64","HU21",2006,5.8,"Közép-Dunántúl"
"Y20-64","HU22",2006,5.6,"Nyugat-Dunántúl"
"Y20-64","HU23",2006,9,"Dél-Dunántúl"
"Y20-64","HU3",2006,9.7,"Alföld és Észak"
"Y20-64","HU31",2006,10.5,"Észak-Magyarország"
"Y20-64","HU32",2006,10.6,"Észak-Alföld"
"Y20-64","HU33",2006,7.9,"Dél-Alföld"
"Y20-64","IE",2006,4.1,"Ireland"
"Y20-64","IE0",2006,4.1,"Éire/Ireland"
"Y20-64","IE01",2006,4.3,"Border, Midland and Western"
"Y20-64","IE02",2006,4,"Southern and Eastern"
"Y20-64","IS",2006,2,"Iceland"
"Y20-64","IS0",2006,2,"Ísland"
"Y20-64","IS00",2006,2,"Ísland"
"Y20-64","IT",2006,6.5,"Italy"
"Y20-64","ITC",2006,3.7,"Nord-Ovest"
"Y20-64","ITC1",2006,3.8,"Piemonte"
"Y20-64","ITC2",2006,2.9,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2006,4.8,"Liguria"
"Y20-64","ITC4",2006,3.5,"Lombardia"
"Y20-64","ITF",2006,11.5,"Sud"
"Y20-64","ITF1",2006,6.5,"Abruzzo"
"Y20-64","ITF2",2006,9.5,"Molise"
"Y20-64","ITF3",2006,12.3,"Campania"
"Y20-64","ITF4",2006,12.1,"Puglia"
"Y20-64","ITF5",2006,10.2,"Basilicata"
"Y20-64","ITF6",2006,12.4,"Calabria"
"Y20-64","ITG",2006,12.1,"Isole"
"Y20-64","ITG1",2006,12.7,"Sicilia"
"Y20-64","ITG2",2006,10.4,"Sardegna"
"Y20-64","ITH",2006,3.4,"Nord-Est"
"Y20-64","ITH1",2006,2.5,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2006,2.9,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2006,3.9,"Veneto"
"Y20-64","ITH4",2006,3.1,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2006,3.2,"Emilia-Romagna"
"Y20-64","ITI",2006,5.9,"Centro (IT)"
"Y20-64","ITI1",2006,4.5,"Toscana"
"Y20-64","ITI2",2006,5,"Umbria"
"Y20-64","ITI3",2006,4.5,"Marche"
"Y20-64","ITI4",2006,7.3,"Lazio"
"Y20-64","LT",2006,5.7,"Lithuania"
"Y20-64","LT0",2006,5.7,"Lietuva"
"Y20-64","LT00",2006,5.7,"Lietuva"
"Y20-64","LU",2006,4.4,"Luxembourg"
"Y20-64","LU0",2006,4.4,"Luxembourg"
"Y20-64","LU00",2006,4.4,"Luxembourg"
"Y20-64","LV",2006,6.7,"Latvia"
"Y20-64","LV0",2006,6.7,"Latvija"
"Y20-64","LV00",2006,6.7,"Latvija"
"Y20-64","MK",2006,35.4,"Former Yugoslav Republic of Macedonia, the"
"Y20-64","MK0",2006,35.4,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MK00",2006,35.4,"Poranesna jugoslovenska Republika Makedonija"
"Y20-64","MT",2006,5.6,"Malta"
"Y20-64","MT0",2006,5.6,"Malta"
"Y20-64","MT00",2006,5.6,"Malta"
"Y20-64","NL",2006,3.5,"Netherlands"
"Y20-64","NL1",2006,4.1,"Noord-Nederland"
"Y20-64","NL11",2006,4.6,"Groningen"
"Y20-64","NL12",2006,3.8,"Friesland (NL)"
"Y20-64","NL13",2006,4,"Drenthe"
"Y20-64","NL2",2006,3.4,"Oost-Nederland"
"Y20-64","NL21",2006,3.7,"Overijssel"
"Y20-64","NL22",2006,3,"Gelderland"
"Y20-64","NL23",2006,4.5,"Flevoland"
"Y20-64","NL3",2006,3.5,"West-Nederland"
"Y20-64","NL31",2006,2.8,"Utrecht"
"Y20-64","NL32",2006,3.4,"Noord-Holland"
"Y20-64","NL33",2006,4,"Zuid-Holland"
"Y20-64","NL34",2006,2.4,"Zeeland"
"Y20-64","NL4",2006,3.4,"Zuid-Nederland"
"Y20-64","NL41",2006,3.1,"Noord-Brabant"
"Y20-64","NL42",2006,4.2,"Limburg (NL)"
"Y20-64","NO",2006,3,"Norway"
"Y20-64","NO0",2006,3,"Norge"
"Y20-64","NO01",2006,3.2,"Oslo og Akershus"
"Y20-64","NO02",2006,2.7,"Hedmark og Oppland"
"Y20-64","NO03",2006,3.4,"Sør-Østlandet"
"Y20-64","NO04",2006,2.5,"Agder og Rogaland"
"Y20-64","NO05",2006,2.4,"Vestlandet"
"Y20-64","NO06",2006,3.1,"Trøndelag"
"Y20-64","NO07",2006,3.2,"Nord-Norge"
"Y20-64","PL",2006,13.8,"Poland"
"Y20-64","PL1",2006,12.6,"Region Centralny"
"Y20-64","PL11",2006,13.5,"Lódzkie"
"Y20-64","PL12",2006,12.2,"Mazowieckie"
"Y20-64","PL2",2006,13.5,"Region Poludniowy"
"Y20-64","PL21",2006,12.7,"Malopolskie"
"Y20-64","PL22",2006,14.1,"Slaskie"
"Y20-64","PL3",2006,13.6,"Region Wschodni"
"Y20-64","PL31",2006,13,"Lubelskie"
"Y20-64","PL32",2006,13.8,"Podkarpackie"
"Y20-64","PL33",2006,15.8,"Swietokrzyskie"
"Y20-64","PL34",2006,11.6,"Podlaskie"
"Y20-64","PL4",2006,13.9,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2006,12.4,"Wielkopolskie"
"Y20-64","PL42",2006,17.1,"Zachodniopomorskie"
"Y20-64","PL43",2006,14,"Lubuskie"
"Y20-64","PL5",2006,16.3,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2006,17.1,"Dolnoslaskie"
"Y20-64","PL52",2006,13.5,"Opolskie"
"Y20-64","PL6",2006,15.1,"Region Pólnocny"
"Y20-64","PL61",2006,16.1,"Kujawsko-Pomorskie"
"Y20-64","PL62",2006,15.7,"Warminsko-Mazurskie"
"Y20-64","PL63",2006,13.6,"Pomorskie"
"Y20-64","PT",2006,7.8,"Portugal"
"Y20-64","PT1",2006,7.9,"Continente"
"Y20-64","PT11",2006,9,"Norte"
"Y20-64","PT15",2006,5.6,"Algarve"
"Y20-64","PT16",2006,6,"Centro (PT)"
"Y20-64","PT17",2006,8.3,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2006,9,"Alentejo"
"Y20-64","PT2",2006,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2006,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2006,5.2,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2006,5.2,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2006,7,"Romania"
"Y20-64","RO1",2006,7.1,"Macroregiunea unu"
"Y20-64","RO11",2006,5.7,"Nord-Vest"
"Y20-64","RO12",2006,8.5,"Centru"
"Y20-64","RO2",2006,7,"Macroregiunea doi"
"Y20-64","RO21",2006,5.9,"Nord-Est"
"Y20-64","RO22",2006,8.6,"Sud-Est"
"Y20-64","RO3",2006,7.1,"Macroregiunea trei"
"Y20-64","RO31",2006,9.1,"Sud - Muntenia"
"Y20-64","RO32",2006,4.5,"Bucuresti - Ilfov"
"Y20-64","RO4",2006,6.9,"Macroregiunea patru"
"Y20-64","RO41",2006,7.5,"Sud-Vest Oltenia"
"Y20-64","RO42",2006,6.2,"Vest"
"Y20-64","SE",2006,6.1,"Sweden"
"Y20-64","SE1",2006,5.7,"Östra Sverige"
"Y20-64","SE11",2006,5.3,"Stockholm"
"Y20-64","SE12",2006,6.4,"Östra Mellansverige"
"Y20-64","SE2",2006,5.9,"Södra Sverige"
"Y20-64","SE21",2006,5,"Småland med öarna"
"Y20-64","SE22",2006,6.9,"Sydsverige"
"Y20-64","SE23",2006,5.7,"Västsverige"
"Y20-64","SE3",2006,7.1,"Norra Sverige"
"Y20-64","SE31",2006,7,"Norra Mellansverige"
"Y20-64","SE32",2006,6.7,"Mellersta Norrland"
"Y20-64","SE33",2006,7.4,"Övre Norrland"
"Y20-64","SI",2006,5.9,"Slovenia"
"Y20-64","SI0",2006,5.9,"Slovenija"
"Y20-64","SI01",2006,7,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2006,4.6,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2006,12.8,"Slovakia"
"Y20-64","SK0",2006,12.8,"Slovensko"
"Y20-64","SK01",2006,4.6,"Bratislavský kraj"
"Y20-64","SK02",2006,9.5,"Západné Slovensko"
"Y20-64","SK03",2006,15.8,"Stredné Slovensko"
"Y20-64","SK04",2006,18.1,"Východné Slovensko"
"Y20-64","TR",2006,8.4,"Turkey"
"Y20-64","TR1",2006,10.1,"Istanbul"
"Y20-64","TR10",2006,10.1,"Istanbul"
"Y20-64","TR2",2006,5.6,"Bati Marmara"
"Y20-64","TR21",2006,6.4,"Tekirdag, Edirne, Kirklareli"
"Y20-64","TR22",2006,4.8,"Balikesir, Çanakkale"
"Y20-64","TR3",2006,7.3,"Ege"
"Y20-64","TR31",2006,9.9,"Izmir"
"Y20-64","TR32",2006,5.1,"Aydin, Denizli, Mugla"
"Y20-64","TR33",2006,6,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y20-64","TR4",2006,8.2,"Dogu Marmara"
"Y20-64","TR41",2006,6.8,"Bursa, Eskisehir, Bilecik"
"Y20-64","TR42",2006,9.9,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y20-64","TR5",2006,10.3,"Bati Anadolu"
"Y20-64","TR51",2006,10.9,"Ankara"
"Y20-64","TR52",2006,8.7,"Konya, Karaman"
"Y20-64","TR6",2006,10.1,"Akdeniz"
"Y20-64","TR61",2006,6.2,"Antalya, Isparta, Burdur"
"Y20-64","TR62",2006,13.9,"Adana, Mersin"
"Y20-64","TR63",2006,9.4,"Hatay, Kahramanmaras, Osmaniye"
"Y20-64","TR7",2006,9,"Orta Anadolu"
"Y20-64","TR71",2006,8.9,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y20-64","TR72",2006,9.1,"Kayseri, Sivas, Yozgat"
"Y20-64","TR8",2006,5.3,"Bati Karadeniz"
"Y20-64","TR81",2006,4.8,"Zonguldak, Karabük, Bartin"
"Y20-64","TR82",2006,3.9,"Kastamonu, Çankiri, Sinop"
"Y20-64","TR83",2006,5.8,"Samsun, Tokat, Çorum, Amasya"
"Y20-64","TR9",2006,4.3,"Dogu Karadeniz"
"Y20-64","TR90",2006,4.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y20-64","TRA",2006,3.5,"Kuzeydogu Anadolu"
"Y20-64","TRA1",2006,3.9,"Erzurum, Erzincan, Bayburt"
"Y20-64","TRA2",2006,3.1,"Agri, Kars, Igdir, Ardahan"
"Y20-64","TRB",2006,8.5,"Ortadogu Anadolu"
"Y20-64","TRB1",2006,10.2,"Malatya, Elazig, Bingöl, Tunceli"
"Y20-64","TRB2",2006,6.6,"Van, Mus, Bitlis, Hakkari"
"Y20-64","TRC",2006,11.8,"Güneydogu Anadolu"
"Y20-64","TRC1",2006,12.6,"Gaziantep, Adiyaman, Kilis"
"Y20-64","TRC2",2006,10.1,"Sanliurfa, Diyarbakir"
"Y20-64","TRC3",2006,13,"Mardin, Batman, Sirnak, Siirt"
"Y20-64","UK",2006,4.5,"United Kingdom"
"Y20-64","UKC",2006,5.3,"North East (UK)"
"Y20-64","UKC1",2006,4.4,"Tees Valley and Durham"
"Y20-64","UKC2",2006,6.1,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2006,4.2,"North West (UK)"
"Y20-64","UKD1",2006,3.5,"Cumbria"
"Y20-64","UKD3",2006,4.5,"Greater Manchester"
"Y20-64","UKD4",2006,4.1,"Lancashire"
"Y20-64","UKD6",2006,2.7,"Cheshire"
"Y20-64","UKD7",2006,5.2,"Merseyside"
"Y20-64","UKE",2006,4.8,"Yorkshire and The Humber"
"Y20-64","UKE1",2006,5,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2006,3.6,"North Yorkshire"
"Y20-64","UKE3",2006,5.7,"South Yorkshire"
"Y20-64","UKE4",2006,4.6,"West Yorkshire"
"Y20-64","UKF",2006,4.2,"East Midlands (UK)"
"Y20-64","UKF1",2006,4.5,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2006,4,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2006,3.6,"Lincolnshire"
"Y20-64","UKG",2006,4.8,"West Midlands (UK)"
"Y20-64","UKG1",2006,3.1,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2006,3.3,"Shropshire and Staffordshire"
"Y20-64","UKG3",2006,6.7,"West Midlands"
"Y20-64","UKH",2006,4,"East of England"
"Y20-64","UKH1",2006,4.1,"East Anglia"
"Y20-64","UKH2",2006,4.2,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2006,3.8,"Essex"
"Y20-64","UKI",2006,6.9,"London"
"Y20-64","UKI1",2006,8.2,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2006,5.9,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2006,3.7,"South East (UK)"
"Y20-64","UKJ1",2006,3.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2006,3.7,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2006,3.9,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2006,4.6,"Kent"
"Y20-64","UKK",2006,3.1,"South West (UK)"
"Y20-64","UKK1",2006,2.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2006,3.2,"Dorset and Somerset"
"Y20-64","UKK3",2006,3.5,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2006,3.5,"Devon"
"Y20-64","UKL",2006,4.3,"Wales"
"Y20-64","UKL1",2006,4.4,"West Wales and The Valleys"
"Y20-64","UKL2",2006,4.2,"East Wales"
"Y20-64","UKM",2006,4.3,"Scotland"
"Y20-64","UKM2",2006,4.2,"Eastern Scotland"
"Y20-64","UKM3",2006,5.1,"South Western Scotland"
"Y20-64","UKM5",2006,1.8,"North Eastern Scotland"
"Y20-64","UKM6",2006,2.9,"Highlands and Islands"
"Y20-64","UKN",2006,3.8,"Northern Ireland (UK)"
"Y20-64","UKN0",2006,3.8,"Northern Ireland (UK)"
"Y_GE15","AT",2006,5.2,"Austria"
"Y_GE15","AT1",2006,7,"Ostösterreich"
"Y_GE15","AT11",2006,5.3,"Burgenland (AT)"
"Y_GE15","AT12",2006,4.5,"Niederösterreich"
"Y_GE15","AT13",2006,9.7,"Wien"
"Y_GE15","AT2",2006,4.4,"Südösterreich"
"Y_GE15","AT21",2006,4.7,"Kärnten"
"Y_GE15","AT22",2006,4.3,"Steiermark"
"Y_GE15","AT3",2006,3.7,"Westösterreich"
"Y_GE15","AT31",2006,3.6,"Oberösterreich"
"Y_GE15","AT32",2006,3.5,"Salzburg"
"Y_GE15","AT33",2006,3.2,"Tirol"
"Y_GE15","AT34",2006,5,"Vorarlberg"
"Y_GE15","BE",2006,8.2,"Belgium"
"Y_GE15","BE1",2006,17.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2006,17.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2006,5,"Vlaams Gewest"
"Y_GE15","BE21",2006,5.7,"Prov. Antwerpen"
"Y_GE15","BE22",2006,6.2,"Prov. Limburg (BE)"
"Y_GE15","BE23",2006,4.5,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2006,4.2,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2006,4.2,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2006,11.7,"Région wallonne"
"Y_GE15","BE31",2006,7.6,"Prov. Brabant Wallon"
"Y_GE15","BE32",2006,14.4,"Prov. Hainaut"
"Y_GE15","BE33",2006,11.5,"Prov. Liège"
"Y_GE15","BE34",2006,7.7,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2006,10.6,"Prov. Namur"
"Y_GE15","BG",2006,9,"Bulgaria"
"Y_GE15","BG3",2006,10.8,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2006,11,"Severozapaden"
"Y_GE15","BG32",2006,13.5,"Severen tsentralen"
"Y_GE15","BG33",2006,11,"Severoiztochen"
"Y_GE15","BG34",2006,8.1,"Yugoiztochen"
"Y_GE15","BG4",2006,7.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2006,6.5,"Yugozapaden"
"Y_GE15","BG42",2006,8.2,"Yuzhen tsentralen"
"Y_GE15","CH",2006,4,"Switzerland"
"Y_GE15","CH0",2006,4,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2006,5.2,"Région lémanique"
"Y_GE15","CH02",2006,3.7,"Espace Mittelland"
"Y_GE15","CH03",2006,4,"Nordwestschweiz"
"Y_GE15","CH04",2006,3.8,"Zürich"
"Y_GE15","CH05",2006,3.6,"Ostschweiz"
"Y_GE15","CH06",2006,2.7,"Zentralschweiz"
"Y_GE15","CH07",2006,5.3,"Ticino"
"Y_GE15","CY",2006,4.5,"Cyprus"
"Y_GE15","CY0",2006,4.5,"Kypros"
"Y_GE15","CY00",2006,4.5,"Kypros"
"Y_GE15","CZ",2006,7.1,"Czech Republic"
"Y_GE15","CZ0",2006,7.1,"Ceská republika"
"Y_GE15","CZ01",2006,2.8,"Praha"
"Y_GE15","CZ02",2006,4.6,"Strední Cechy"
"Y_GE15","CZ03",2006,4.9,"Jihozápad"
"Y_GE15","CZ04",2006,12.8,"Severozápad"
"Y_GE15","CZ05",2006,6.1,"Severovýchod"
"Y_GE15","CZ06",2006,7.1,"Jihovýchod"
"Y_GE15","CZ07",2006,7.6,"Strední Morava"
"Y_GE15","CZ08",2006,12,"Moravskoslezsko"
"Y_GE15","DE",2006,10.3,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2006,6.4,"Baden-Württemberg"
"Y_GE15","DE11",2006,6.5,"Stuttgart"
"Y_GE15","DE12",2006,7.2,"Karlsruhe"
"Y_GE15","DE13",2006,5.5,"Freiburg"
"Y_GE15","DE14",2006,5.9,"Tübingen"
"Y_GE15","DE2",2006,6.5,"Bayern"
"Y_GE15","DE21",2006,5.3,"Oberbayern"
"Y_GE15","DE22",2006,6.6,"Niederbayern"
"Y_GE15","DE23",2006,6.8,"Oberpfalz"
"Y_GE15","DE24",2006,9.6,"Oberfranken"
"Y_GE15","DE25",2006,7.9,"Mittelfranken"
"Y_GE15","DE26",2006,6.3,"Unterfranken"
"Y_GE15","DE27",2006,6.2,"Schwaben"
"Y_GE15","DE3",2006,18.7,"Berlin"
"Y_GE15","DE30",2006,18.7,"Berlin"
"Y_GE15","DE4",2006,16.6,"Brandenburg"
"Y_GE15","DE40",2006,16.6,"Brandenburg"
"Y_GE15","DE5",2006,14.4,"Bremen"
"Y_GE15","DE50",2006,14.4,"Bremen"
"Y_GE15","DE6",2006,9.9,"Hamburg"
"Y_GE15","DE60",2006,9.9,"Hamburg"
"Y_GE15","DE7",2006,8.1,"Hessen"
"Y_GE15","DE71",2006,7.9,"Darmstadt"
"Y_GE15","DE72",2006,8.5,"Gießen"
"Y_GE15","DE73",2006,8.5,"Kassel"
"Y_GE15","DE8",2006,19.2,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2006,19.2,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2006,9.7,"Niedersachsen"
"Y_GE15","DE91",2006,10.1,"Braunschweig"
"Y_GE15","DE92",2006,10.5,"Hannover"
"Y_GE15","DE93",2006,9,"Lüneburg"
"Y_GE15","DE94",2006,9.3,"Weser-Ems"
"Y_GE15","DEA",2006,9.8,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2006,9.8,"Düsseldorf"
"Y_GE15","DEA2",2006,9.1,"Köln"
"Y_GE15","DEA3",2006,9.1,"Münster"
"Y_GE15","DEA4",2006,10,"Detmold"
"Y_GE15","DEA5",2006,11.1,"Arnsberg"
"Y_GE15","DEB",2006,8,"Rheinland-Pfalz"
"Y_GE15","DEB1",2006,7.8,"Koblenz"
"Y_GE15","DEB2",2006,6.2,"Trier"
"Y_GE15","DEB3",2006,8.7,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2006,9.5,"Saarland"
"Y_GE15","DEC0",2006,9.5,"Saarland"
"Y_GE15","DED",2006,16.7,"Sachsen"
"Y_GE15","DED2",2006,16.2,"Dresden"
"Y_GE15","DED4",2006,16.5,"Chemnitz"
"Y_GE15","DED5",2006,17.8,"Leipzig"
"Y_GE15","DEE",2006,17.8,"Sachsen-Anhalt"
"Y_GE15","DEE0",2006,17.8,"Sachsen-Anhalt"
"Y_GE15","DEF",2006,9.1,"Schleswig-Holstein"
"Y_GE15","DEF0",2006,9.1,"Schleswig-Holstein"
"Y_GE15","DEG",2006,15.7,"Thüringen"
"Y_GE15","DEG0",2006,15.7,"Thüringen"
"Y_GE15","DK",2006,3.9,"Denmark"
"Y_GE15","DK0",2006,3.9,"Danmark"
"Y_GE15","EA17",2006,8.4,"Euro area (17 countries)"
"Y_GE15","EA18",2006,8.4,"Euro area (18 countries)"
"Y_GE15","EA19",2006,8.3,"Euro area (19 countries)"
"Y_GE15","EE",2006,5.9,"Estonia"
"Y_GE15","EE0",2006,5.9,"Eesti"
"Y_GE15","EE00",2006,5.9,"Eesti"
"Y_GE15","EL",2006,9,"Greece"
"Y_GE15","EL1",2006,9.8,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2006,11.1,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2006,9.5,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2006,14.2,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2006,8.2,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2006,9.2,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2006,9.8,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2006,11.2,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2006,9.7,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2006,9.2,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2006,7.5,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2006,8.5,"Attiki"
"Y_GE15","EL30",2006,8.5,"Attiki"
"Y_GE15","EL4",2006,8.1,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2006,9.6,"Voreio Aigaio"
"Y_GE15","EL42",2006,9,"Notio Aigaio"
"Y_GE15","EL43",2006,7.2,"Kriti"
"Y_GE15","ES",2006,8.5,"Spain"
"Y_GE15","ES1",2006,8.3,"Noroeste (ES)"
"Y_GE15","ES11",2006,8.3,"Galicia"
"Y_GE15","ES12",2006,9.2,"Principado de Asturias"
"Y_GE15","ES13",2006,6.5,"Cantabria"
"Y_GE15","ES2",2006,6.4,"Noreste (ES)"
"Y_GE15","ES21",2006,7.2,"País Vasco"
"Y_GE15","ES22",2006,5.4,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2006,6.1,"La Rioja"
"Y_GE15","ES24",2006,5.5,"Aragón"
"Y_GE15","ES3",2006,6.3,"Comunidad de Madrid"
"Y_GE15","ES30",2006,6.3,"Comunidad de Madrid"
"Y_GE15","ES4",2006,9.3,"Centro (ES)"
"Y_GE15","ES41",2006,8.1,"Castilla y León"
"Y_GE15","ES42",2006,8.8,"Castilla-la Mancha"
"Y_GE15","ES43",2006,13.3,"Extremadura"
"Y_GE15","ES5",2006,7.1,"Este (ES)"
"Y_GE15","ES51",2006,6.5,"Cataluña"
"Y_GE15","ES52",2006,8.3,"Comunidad Valenciana"
"Y_GE15","ES53",2006,6.4,"Illes Balears"
"Y_GE15","ES6",2006,12,"Sur (ES)"
"Y_GE15","ES61",2006,12.6,"Andalucía"
"Y_GE15","ES62",2006,7.9,"Región de Murcia"
"Y_GE15","ES63",2006,21.5,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2006,13.6,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2006,11.6,"Canarias (ES)"
"Y_GE15","ES70",2006,11.6,"Canarias (ES)"
"Y_GE15","EU15",2006,7.7,"European Union (15 countries)"
"Y_GE15","EU27",2006,8.2,"European Union (27 countries)"
"Y_GE15","EU28",2006,8.2,"European Union (28 countries)"
"Y_GE15","FI",2006,7.7,"Finland"
"Y_GE15","FI1",2006,7.7,"Manner-Suomi"
"Y_GE15","FI19",2006,7.8,"Länsi-Suomi"
"Y_GE15","FI1B",2006,5.4,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2006,7.7,"Etelä-Suomi"
"Y_GE15","FI1D",2006,10.8,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2006,NA,"Åland"
"Y_GE15","FI20",2006,NA,"Åland"
"Y_GE15","FR",2006,8.9,"France"
"Y_GE15","FR1",2006,8.5,"Île de France"
"Y_GE15","FR10",2006,8.5,"Île de France"
"Y_GE15","FR2",2006,8.1,"Bassin Parisien"
"Y_GE15","FR21",2006,6.8,"Champagne-Ardenne"
"Y_GE15","FR22",2006,10.2,"Picardie"
"Y_GE15","FR23",2006,8.8,"Haute-Normandie"
"Y_GE15","FR24",2006,6.9,"Centre (FR)"
"Y_GE15","FR25",2006,7.2,"Basse-Normandie"
"Y_GE15","FR26",2006,8.4,"Bourgogne"
"Y_GE15","FR3",2006,12,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2006,12,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2006,8,"Est (FR)"
"Y_GE15","FR41",2006,9.5,"Lorraine"
"Y_GE15","FR42",2006,6.4,"Alsace"
"Y_GE15","FR43",2006,7.6,"Franche-Comté"
"Y_GE15","FR5",2006,7.2,"Ouest (FR)"
"Y_GE15","FR51",2006,6.9,"Pays de la Loire"
"Y_GE15","FR52",2006,7.3,"Bretagne"
"Y_GE15","FR53",2006,7.7,"Poitou-Charentes"
"Y_GE15","FR6",2006,7.5,"Sud-Ouest (FR)"
"Y_GE15","FR61",2006,7.5,"Aquitaine"
"Y_GE15","FR62",2006,7.9,"Midi-Pyrénées"
"Y_GE15","FR63",2006,5.8,"Limousin"
"Y_GE15","FR7",2006,7.3,"Centre-Est (FR)"
"Y_GE15","FR71",2006,7.3,"Rhône-Alpes"
"Y_GE15","FR72",2006,7.3,"Auvergne"
"Y_GE15","FR8",2006,11,"Méditerranée"
"Y_GE15","FR81",2006,10.9,"Languedoc-Roussillon"
"Y_GE15","FR82",2006,11,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2006,10.7,"Corse"
"Y_GE15","FR9",2006,27,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2006,26.9,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2006,24.1,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2006,28.5,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2006,28.3,"Réunion (NUTS 2010)"
"Y_GE15","HR",2006,11.1,"Croatia"
"Y_GE15","HR0",2006,11.1,"Hrvatska"
"Y_GE15","HU",2006,7.5,"Hungary"
"Y_GE15","HU1",2006,5.1,"Közép-Magyarország"
"Y_GE15","HU10",2006,5.1,"Közép-Magyarország"
"Y_GE15","HU2",2006,6.9,"Dunántúl"
"Y_GE15","HU21",2006,6,"Közép-Dunántúl"
"Y_GE15","HU22",2006,5.8,"Nyugat-Dunántúl"
"Y_GE15","HU23",2006,9.2,"Dél-Dunántúl"
"Y_GE15","HU3",2006,10,"Alföld és Észak"
"Y_GE15","HU31",2006,10.9,"Észak-Magyarország"
"Y_GE15","HU32",2006,10.9,"Észak-Alföld"
"Y_GE15","HU33",2006,8,"Dél-Alföld"
"Y_GE15","IE",2006,4.4,"Ireland"
"Y_GE15","IE0",2006,4.4,"Éire/Ireland"
"Y_GE15","IE01",2006,4.7,"Border, Midland and Western"
"Y_GE15","IE02",2006,4.3,"Southern and Eastern"
"Y_GE15","IS",2006,2.8,"Iceland"
"Y_GE15","IS0",2006,2.8,"Ísland"
"Y_GE15","IS00",2006,2.8,"Ísland"
"Y_GE15","IT",2006,6.8,"Italy"
"Y_GE15","ITC",2006,3.9,"Nord-Ovest"
"Y_GE15","ITC1",2006,4.1,"Piemonte"
"Y_GE15","ITC2",2006,2.9,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2006,4.8,"Liguria"
"Y_GE15","ITC4",2006,3.7,"Lombardia"
"Y_GE15","ITF",2006,11.9,"Sud"
"Y_GE15","ITF1",2006,6.6,"Abruzzo"
"Y_GE15","ITF2",2006,9.9,"Molise"
"Y_GE15","ITF3",2006,12.8,"Campania"
"Y_GE15","ITF4",2006,12.6,"Puglia"
"Y_GE15","ITF5",2006,10.6,"Basilicata"
"Y_GE15","ITF6",2006,12.8,"Calabria"
"Y_GE15","ITG",2006,12.7,"Isole"
"Y_GE15","ITG1",2006,13.4,"Sicilia"
"Y_GE15","ITG2",2006,10.7,"Sardegna"
"Y_GE15","ITH",2006,3.6,"Nord-Est"
"Y_GE15","ITH1",2006,2.6,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2006,3.1,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2006,4.1,"Veneto"
"Y_GE15","ITH4",2006,3.5,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2006,3.4,"Emilia-Romagna"
"Y_GE15","ITI",2006,6.1,"Centro (IT)"
"Y_GE15","ITI1",2006,4.8,"Toscana"
"Y_GE15","ITI2",2006,5.1,"Umbria"
"Y_GE15","ITI3",2006,4.6,"Marche"
"Y_GE15","ITI4",2006,7.5,"Lazio"
"Y_GE15","LT",2006,5.8,"Lithuania"
"Y_GE15","LT0",2006,5.8,"Lietuva"
"Y_GE15","LT00",2006,5.8,"Lietuva"
"Y_GE15","LU",2006,4.7,"Luxembourg"
"Y_GE15","LU0",2006,4.7,"Luxembourg"
"Y_GE15","LU00",2006,4.7,"Luxembourg"
"Y_GE15","LV",2006,7,"Latvia"
"Y_GE15","LV0",2006,7,"Latvija"
"Y_GE15","LV00",2006,7,"Latvija"
"Y_GE15","MK",2006,36,"Former Yugoslav Republic of Macedonia, the"
"Y_GE15","MK0",2006,36,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MK00",2006,36,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE15","MT",2006,6.8,"Malta"
"Y_GE15","MT0",2006,6.8,"Malta"
"Y_GE15","MT00",2006,6.8,"Malta"
"Y_GE15","NL",2006,3.9,"Netherlands"
"Y_GE15","NL1",2006,4.6,"Noord-Nederland"
"Y_GE15","NL11",2006,5,"Groningen"
"Y_GE15","NL12",2006,4.2,"Friesland (NL)"
"Y_GE15","NL13",2006,4.6,"Drenthe"
"Y_GE15","NL2",2006,3.7,"Oost-Nederland"
"Y_GE15","NL21",2006,4,"Overijssel"
"Y_GE15","NL22",2006,3.3,"Gelderland"
"Y_GE15","NL23",2006,5.2,"Flevoland"
"Y_GE15","NL3",2006,3.9,"West-Nederland"
"Y_GE15","NL31",2006,3.3,"Utrecht"
"Y_GE15","NL32",2006,3.8,"Noord-Holland"
"Y_GE15","NL33",2006,4.4,"Zuid-Holland"
"Y_GE15","NL34",2006,2.7,"Zeeland"
"Y_GE15","NL4",2006,3.7,"Zuid-Nederland"
"Y_GE15","NL41",2006,3.4,"Noord-Brabant"
"Y_GE15","NL42",2006,4.5,"Limburg (NL)"
"Y_GE15","NO",2006,3.4,"Norway"
"Y_GE15","NO0",2006,3.4,"Norge"
"Y_GE15","NO01",2006,3.5,"Oslo og Akershus"
"Y_GE15","NO02",2006,3.1,"Hedmark og Oppland"
"Y_GE15","NO03",2006,4,"Sør-Østlandet"
"Y_GE15","NO04",2006,2.9,"Agder og Rogaland"
"Y_GE15","NO05",2006,2.8,"Vestlandet"
"Y_GE15","NO06",2006,3.6,"Trøndelag"
"Y_GE15","NO07",2006,3.8,"Nord-Norge"
"Y_GE15","PL",2006,13.8,"Poland"
"Y_GE15","PL1",2006,12.7,"Region Centralny"
"Y_GE15","PL11",2006,13.4,"Lódzkie"
"Y_GE15","PL12",2006,12.3,"Mazowieckie"
"Y_GE15","PL2",2006,13.5,"Region Poludniowy"
"Y_GE15","PL21",2006,12.6,"Malopolskie"
"Y_GE15","PL22",2006,14.2,"Slaskie"
"Y_GE15","PL3",2006,13.4,"Region Wschodni"
"Y_GE15","PL31",2006,12.8,"Lubelskie"
"Y_GE15","PL32",2006,13.7,"Podkarpackie"
"Y_GE15","PL33",2006,15.5,"Swietokrzyskie"
"Y_GE15","PL34",2006,11.3,"Podlaskie"
"Y_GE15","PL4",2006,14.1,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2006,12.7,"Wielkopolskie"
"Y_GE15","PL42",2006,17.2,"Zachodniopomorskie"
"Y_GE15","PL43",2006,14,"Lubuskie"
"Y_GE15","PL5",2006,16.4,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2006,17.3,"Dolnoslaskie"
"Y_GE15","PL52",2006,13.5,"Opolskie"
"Y_GE15","PL6",2006,15.3,"Region Pólnocny"
"Y_GE15","PL61",2006,16.2,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2006,16,"Warminsko-Mazurskie"
"Y_GE15","PL63",2006,13.8,"Pomorskie"
"Y_GE15","PT",2006,7.6,"Portugal"
"Y_GE15","PT1",2006,7.8,"Continente"
"Y_GE15","PT11",2006,8.8,"Norte"
"Y_GE15","PT15",2006,5.5,"Algarve"
"Y_GE15","PT16",2006,5.4,"Centro (PT)"
"Y_GE15","PT17",2006,8.5,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2006,9.1,"Alentejo"
"Y_GE15","PT2",2006,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2006,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2006,5.3,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2006,5.3,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2006,7.3,"Romania"
"Y_GE15","RO1",2006,7.4,"Macroregiunea unu"
"Y_GE15","RO11",2006,5.9,"Nord-Vest"
"Y_GE15","RO12",2006,9,"Centru"
"Y_GE15","RO2",2006,7.2,"Macroregiunea doi"
"Y_GE15","RO21",2006,5.9,"Nord-Est"
"Y_GE15","RO22",2006,9,"Sud-Est"
"Y_GE15","RO3",2006,7.5,"Macroregiunea trei"
"Y_GE15","RO31",2006,9.4,"Sud - Muntenia"
"Y_GE15","RO32",2006,4.8,"Bucuresti - Ilfov"
"Y_GE15","RO4",2006,6.8,"Macroregiunea patru"
"Y_GE15","RO41",2006,7.1,"Sud-Vest Oltenia"
"Y_GE15","RO42",2006,6.4,"Vest"
"Y_GE15","SE",2006,7.1,"Sweden"
"Y_GE15","SE1",2006,6.6,"Östra Sverige"
"Y_GE15","SE11",2006,6.1,"Stockholm"
"Y_GE15","SE12",2006,7.3,"Östra Mellansverige"
"Y_GE15","SE2",2006,7.1,"Södra Sverige"
"Y_GE15","SE21",2006,5.9,"Småland med öarna"
"Y_GE15","SE22",2006,8.2,"Sydsverige"
"Y_GE15","SE23",2006,6.8,"Västsverige"
"Y_GE15","SE3",2006,8,"Norra Sverige"
"Y_GE15","SE31",2006,7.9,"Norra Mellansverige"
"Y_GE15","SE32",2006,7.3,"Mellersta Norrland"
"Y_GE15","SE33",2006,8.5,"Övre Norrland"
"Y_GE15","SI",2006,6,"Slovenia"
"Y_GE15","SI0",2006,6,"Slovenija"
"Y_GE15","SI01",2006,7.1,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2006,4.6,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2006,13.4,"Slovakia"
"Y_GE15","SK0",2006,13.4,"Slovensko"
"Y_GE15","SK01",2006,4.6,"Bratislavský kraj"
"Y_GE15","SK02",2006,9.8,"Západné Slovensko"
"Y_GE15","SK03",2006,16.4,"Stredné Slovensko"
"Y_GE15","SK04",2006,19.1,"Východné Slovensko"
"Y_GE15","TR",2006,8.7,"Turkey"
"Y_GE15","TR1",2006,10.5,"Istanbul"
"Y_GE15","TR10",2006,10.5,"Istanbul"
"Y_GE15","TR2",2006,5.9,"Bati Marmara"
"Y_GE15","TR21",2006,6.8,"Tekirdag, Edirne, Kirklareli"
"Y_GE15","TR22",2006,4.9,"Balikesir, Çanakkale"
"Y_GE15","TR3",2006,7.5,"Ege"
"Y_GE15","TR31",2006,10.3,"Izmir"
"Y_GE15","TR32",2006,5.3,"Aydin, Denizli, Mugla"
"Y_GE15","TR33",2006,6.2,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE15","TR4",2006,8.6,"Dogu Marmara"
"Y_GE15","TR41",2006,7.3,"Bursa, Eskisehir, Bilecik"
"Y_GE15","TR42",2006,10.3,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE15","TR5",2006,10.8,"Bati Anadolu"
"Y_GE15","TR51",2006,11.4,"Ankara"
"Y_GE15","TR52",2006,9.2,"Konya, Karaman"
"Y_GE15","TR6",2006,10.4,"Akdeniz"
"Y_GE15","TR61",2006,6.4,"Antalya, Isparta, Burdur"
"Y_GE15","TR62",2006,14.3,"Adana, Mersin"
"Y_GE15","TR63",2006,9.5,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE15","TR7",2006,9.4,"Orta Anadolu"
"Y_GE15","TR71",2006,9.2,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE15","TR72",2006,9.5,"Kayseri, Sivas, Yozgat"
"Y_GE15","TR8",2006,5.2,"Bati Karadeniz"
"Y_GE15","TR81",2006,4.8,"Zonguldak, Karabük, Bartin"
"Y_GE15","TR82",2006,3.9,"Kastamonu, Çankiri, Sinop"
"Y_GE15","TR83",2006,5.7,"Samsun, Tokat, Çorum, Amasya"
"Y_GE15","TR9",2006,4.3,"Dogu Karadeniz"
"Y_GE15","TR90",2006,4.3,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE15","TRA",2006,3.6,"Kuzeydogu Anadolu"
"Y_GE15","TRA1",2006,3.9,"Erzurum, Erzincan, Bayburt"
"Y_GE15","TRA2",2006,3.3,"Agri, Kars, Igdir, Ardahan"
"Y_GE15","TRB",2006,8.8,"Ortadogu Anadolu"
"Y_GE15","TRB1",2006,10.5,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE15","TRB2",2006,6.9,"Van, Mus, Bitlis, Hakkari"
"Y_GE15","TRC",2006,12.1,"Güneydogu Anadolu"
"Y_GE15","TRC1",2006,12.6,"Gaziantep, Adiyaman, Kilis"
"Y_GE15","TRC2",2006,10.8,"Sanliurfa, Diyarbakir"
"Y_GE15","TRC3",2006,13.5,"Mardin, Batman, Sirnak, Siirt"
"Y_GE15","UK",2006,5.3,"United Kingdom"
"Y_GE15","UKC",2006,6.4,"North East (UK)"
"Y_GE15","UKC1",2006,5.8,"Tees Valley and Durham"
"Y_GE15","UKC2",2006,6.9,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2006,5.1,"North West (UK)"
"Y_GE15","UKD1",2006,4.3,"Cumbria"
"Y_GE15","UKD3",2006,5.4,"Greater Manchester"
"Y_GE15","UKD4",2006,4.9,"Lancashire"
"Y_GE15","UKD6",2006,3.3,"Cheshire"
"Y_GE15","UKD7",2006,6.4,"Merseyside"
"Y_GE15","UKE",2006,5.7,"Yorkshire and The Humber"
"Y_GE15","UKE1",2006,6,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2006,4,"North Yorkshire"
"Y_GE15","UKE3",2006,7,"South Yorkshire"
"Y_GE15","UKE4",2006,5.5,"West Yorkshire"
"Y_GE15","UKF",2006,5.2,"East Midlands (UK)"
"Y_GE15","UKF1",2006,5.5,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2006,5.1,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2006,4.7,"Lincolnshire"
"Y_GE15","UKG",2006,5.8,"West Midlands (UK)"
"Y_GE15","UKG1",2006,3.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2006,4.2,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2006,7.9,"West Midlands"
"Y_GE15","UKH",2006,4.7,"East of England"
"Y_GE15","UKH1",2006,4.7,"East Anglia"
"Y_GE15","UKH2",2006,4.8,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2006,4.6,"Essex"
"Y_GE15","UKI",2006,7.8,"London"
"Y_GE15","UKI1",2006,8.8,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2006,7.1,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2006,4.4,"South East (UK)"
"Y_GE15","UKJ1",2006,3.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2006,4,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2006,4.6,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2006,5.5,"Kent"
"Y_GE15","UKK",2006,3.7,"South West (UK)"
"Y_GE15","UKK1",2006,3.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2006,3.7,"Dorset and Somerset"
"Y_GE15","UKK3",2006,3.9,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2006,4.4,"Devon"
"Y_GE15","UKL",2006,5.2,"Wales"
"Y_GE15","UKL1",2006,5.4,"West Wales and The Valleys"
"Y_GE15","UKL2",2006,4.9,"East Wales"
"Y_GE15","UKM",2006,5.2,"Scotland"
"Y_GE15","UKM2",2006,5.3,"Eastern Scotland"
"Y_GE15","UKM3",2006,6,"South Western Scotland"
"Y_GE15","UKM5",2006,2.6,"North Eastern Scotland"
"Y_GE15","UKM6",2006,3.2,"Highlands and Islands"
"Y_GE15","UKN",2006,4.3,"Northern Ireland (UK)"
"Y_GE15","UKN0",2006,4.3,"Northern Ireland (UK)"
"Y_GE25","AT",2006,4.5,"Austria"
"Y_GE25","AT1",2006,6,"Ostösterreich"
"Y_GE25","AT11",2006,4.4,"Burgenland (AT)"
"Y_GE25","AT12",2006,3.8,"Niederösterreich"
"Y_GE25","AT13",2006,8.4,"Wien"
"Y_GE25","AT2",2006,3.8,"Südösterreich"
"Y_GE25","AT21",2006,4.1,"Kärnten"
"Y_GE25","AT22",2006,3.7,"Steiermark"
"Y_GE25","AT3",2006,3.1,"Westösterreich"
"Y_GE25","AT31",2006,3.1,"Oberösterreich"
"Y_GE25","AT32",2006,2.9,"Salzburg"
"Y_GE25","AT33",2006,2.6,"Tirol"
"Y_GE25","AT34",2006,4.3,"Vorarlberg"
"Y_GE25","BE",2006,7,"Belgium"
"Y_GE25","BE1",2006,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2006,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2006,4.2,"Vlaams Gewest"
"Y_GE25","BE21",2006,4.9,"Prov. Antwerpen"
"Y_GE25","BE22",2006,5.4,"Prov. Limburg (BE)"
"Y_GE25","BE23",2006,3.9,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2006,3.3,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2006,3.4,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2006,9.6,"Région wallonne"
"Y_GE25","BE31",2006,6.1,"Prov. Brabant Wallon"
"Y_GE25","BE32",2006,11.9,"Prov. Hainaut"
"Y_GE25","BE33",2006,9.5,"Prov. Liège"
"Y_GE25","BE34",2006,5.7,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2006,8.5,"Prov. Namur"
"Y_GE25","BG",2006,7.9,"Bulgaria"
"Y_GE25","BG3",2006,9.6,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2006,9.8,"Severozapaden"
"Y_GE25","BG32",2006,12.2,"Severen tsentralen"
"Y_GE25","BG33",2006,9.7,"Severoiztochen"
"Y_GE25","BG34",2006,7.1,"Yugoiztochen"
"Y_GE25","BG4",2006,6.3,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2006,5.8,"Yugozapaden"
"Y_GE25","BG42",2006,7.1,"Yuzhen tsentralen"
"Y_GE25","CH",2006,3.4,"Switzerland"
"Y_GE25","CH0",2006,3.4,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2006,4.5,"Région lémanique"
"Y_GE25","CH02",2006,3.2,"Espace Mittelland"
"Y_GE25","CH03",2006,3.3,"Nordwestschweiz"
"Y_GE25","CH04",2006,3.1,"Zürich"
"Y_GE25","CH05",2006,2.9,"Ostschweiz"
"Y_GE25","CH06",2006,2.5,"Zentralschweiz"
"Y_GE25","CH07",2006,4.4,"Ticino"
"Y_GE25","CY",2006,3.9,"Cyprus"
"Y_GE25","CY0",2006,3.9,"Kypros"
"Y_GE25","CY00",2006,3.9,"Kypros"
"Y_GE25","CZ",2006,6.2,"Czech Republic"
"Y_GE25","CZ0",2006,6.2,"Ceská republika"
"Y_GE25","CZ01",2006,2.5,"Praha"
"Y_GE25","CZ02",2006,4,"Strední Cechy"
"Y_GE25","CZ03",2006,4.2,"Jihozápad"
"Y_GE25","CZ04",2006,11,"Severozápad"
"Y_GE25","CZ05",2006,5.5,"Severovýchod"
"Y_GE25","CZ06",2006,6,"Jihovýchod"
"Y_GE25","CZ07",2006,6.9,"Strední Morava"
"Y_GE25","CZ08",2006,10,"Moravskoslezsko"
"Y_GE25","DE",2006,9.8,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2006,6,"Baden-Württemberg"
"Y_GE25","DE11",2006,6.1,"Stuttgart"
"Y_GE25","DE12",2006,6.8,"Karlsruhe"
"Y_GE25","DE13",2006,5.4,"Freiburg"
"Y_GE25","DE14",2006,5.4,"Tübingen"
"Y_GE25","DE2",2006,6.2,"Bayern"
"Y_GE25","DE21",2006,5.1,"Oberbayern"
"Y_GE25","DE22",2006,5.8,"Niederbayern"
"Y_GE25","DE23",2006,6.8,"Oberpfalz"
"Y_GE25","DE24",2006,9.2,"Oberfranken"
"Y_GE25","DE25",2006,7.7,"Mittelfranken"
"Y_GE25","DE26",2006,5.7,"Unterfranken"
"Y_GE25","DE27",2006,6,"Schwaben"
"Y_GE25","DE3",2006,18,"Berlin"
"Y_GE25","DE30",2006,18,"Berlin"
"Y_GE25","DE4",2006,16.1,"Brandenburg"
"Y_GE25","DE40",2006,16.1,"Brandenburg"
"Y_GE25","DE5",2006,14.2,"Bremen"
"Y_GE25","DE50",2006,14.2,"Bremen"
"Y_GE25","DE6",2006,9.2,"Hamburg"
"Y_GE25","DE60",2006,9.2,"Hamburg"
"Y_GE25","DE7",2006,7.5,"Hessen"
"Y_GE25","DE71",2006,7.4,"Darmstadt"
"Y_GE25","DE72",2006,7.5,"Gießen"
"Y_GE25","DE73",2006,7.9,"Kassel"
"Y_GE25","DE8",2006,19,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2006,19,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2006,9.2,"Niedersachsen"
"Y_GE25","DE91",2006,9.6,"Braunschweig"
"Y_GE25","DE92",2006,10.2,"Hannover"
"Y_GE25","DE93",2006,8.1,"Lüneburg"
"Y_GE25","DE94",2006,8.9,"Weser-Ems"
"Y_GE25","DEA",2006,9.3,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2006,9.2,"Düsseldorf"
"Y_GE25","DEA2",2006,8.7,"Köln"
"Y_GE25","DEA3",2006,8.3,"Münster"
"Y_GE25","DEA4",2006,9.5,"Detmold"
"Y_GE25","DEA5",2006,10.7,"Arnsberg"
"Y_GE25","DEB",2006,7.3,"Rheinland-Pfalz"
"Y_GE25","DEB1",2006,7.1,"Koblenz"
"Y_GE25","DEB2",2006,5.8,"Trier"
"Y_GE25","DEB3",2006,7.8,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2006,9,"Saarland"
"Y_GE25","DEC0",2006,9,"Saarland"
"Y_GE25","DED",2006,16.5,"Sachsen"
"Y_GE25","DED2",2006,15.8,"Dresden"
"Y_GE25","DED4",2006,16.5,"Chemnitz"
"Y_GE25","DED5",2006,17.6,"Leipzig"
"Y_GE25","DEE",2006,17.7,"Sachsen-Anhalt"
"Y_GE25","DEE0",2006,17.7,"Sachsen-Anhalt"
"Y_GE25","DEF",2006,8.5,"Schleswig-Holstein"
"Y_GE25","DEF0",2006,8.5,"Schleswig-Holstein"
"Y_GE25","DEG",2006,15.4,"Thüringen"
"Y_GE25","DEG0",2006,15.4,"Thüringen"
"Y_GE25","DK",2006,3.2,"Denmark"
"Y_GE25","DK0",2006,3.2,"Danmark"
"Y_GE25","EA17",2006,7.3,"Euro area (17 countries)"
"Y_GE25","EA18",2006,7.3,"Euro area (18 countries)"
"Y_GE25","EA19",2006,7.3,"Euro area (19 countries)"
"Y_GE25","EE",2006,5.2,"Estonia"
"Y_GE25","EE0",2006,5.2,"Eesti"
"Y_GE25","EE00",2006,5.2,"Eesti"
"Y_GE25","EL",2006,7.5,"Greece"
"Y_GE25","EL1",2006,8.2,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2006,8.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2006,7.9,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2006,13.1,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2006,6.7,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2006,7.2,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2006,7.9,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2006,9.2,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2006,7.3,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2006,7.3,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2006,6,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2006,7.3,"Attiki"
"Y_GE25","EL30",2006,7.3,"Attiki"
"Y_GE25","EL4",2006,6.8,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2006,6.9,"Voreio Aigaio"
"Y_GE25","EL42",2006,8,"Notio Aigaio"
"Y_GE25","EL43",2006,6.1,"Kriti"
"Y_GE25","ES",2006,7.2,"Spain"
"Y_GE25","ES1",2006,7.2,"Noroeste (ES)"
"Y_GE25","ES11",2006,7.4,"Galicia"
"Y_GE25","ES12",2006,7.9,"Principado de Asturias"
"Y_GE25","ES13",2006,5.4,"Cantabria"
"Y_GE25","ES2",2006,5.3,"Noreste (ES)"
"Y_GE25","ES21",2006,5.9,"País Vasco"
"Y_GE25","ES22",2006,4.4,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2006,5.1,"La Rioja"
"Y_GE25","ES24",2006,4.8,"Aragón"
"Y_GE25","ES3",2006,5.3,"Comunidad de Madrid"
"Y_GE25","ES30",2006,5.3,"Comunidad de Madrid"
"Y_GE25","ES4",2006,8.1,"Centro (ES)"
"Y_GE25","ES41",2006,7.2,"Castilla y León"
"Y_GE25","ES42",2006,7.6,"Castilla-la Mancha"
"Y_GE25","ES43",2006,11.7,"Extremadura"
"Y_GE25","ES5",2006,6,"Este (ES)"
"Y_GE25","ES51",2006,5.5,"Cataluña"
"Y_GE25","ES52",2006,7,"Comunidad Valenciana"
"Y_GE25","ES53",2006,5.5,"Illes Balears"
"Y_GE25","ES6",2006,10.5,"Sur (ES)"
"Y_GE25","ES61",2006,11.2,"Andalucía"
"Y_GE25","ES62",2006,6.4,"Región de Murcia"
"Y_GE25","ES63",2006,16.1,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2006,11.5,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2006,10,"Canarias (ES)"
"Y_GE25","ES70",2006,10,"Canarias (ES)"
"Y_GE25","EU15",2006,6.6,"European Union (15 countries)"
"Y_GE25","EU27",2006,7,"European Union (27 countries)"
"Y_GE25","EU28",2006,7,"European Union (28 countries)"
"Y_GE25","FI",2006,6.2,"Finland"
"Y_GE25","FI1",2006,6.2,"Manner-Suomi"
"Y_GE25","FI19",2006,6.2,"Länsi-Suomi"
"Y_GE25","FI1B",2006,4.2,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2006,6.4,"Etelä-Suomi"
"Y_GE25","FI1D",2006,8.6,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2006,NA,"Åland"
"Y_GE25","FI20",2006,NA,"Åland"
"Y_GE25","FR",2006,7.3,"France"
"Y_GE25","FR1",2006,7.3,"Île de France"
"Y_GE25","FR10",2006,7.3,"Île de France"
"Y_GE25","FR2",2006,6.4,"Bassin Parisien"
"Y_GE25","FR21",2006,5.4,"Champagne-Ardenne"
"Y_GE25","FR22",2006,8,"Picardie"
"Y_GE25","FR23",2006,6.5,"Haute-Normandie"
"Y_GE25","FR24",2006,5.5,"Centre (FR)"
"Y_GE25","FR25",2006,5.7,"Basse-Normandie"
"Y_GE25","FR26",2006,7.1,"Bourgogne"
"Y_GE25","FR3",2006,9.6,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2006,9.6,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2006,6.2,"Est (FR)"
"Y_GE25","FR41",2006,7.1,"Lorraine"
"Y_GE25","FR42",2006,5.2,"Alsace"
"Y_GE25","FR43",2006,6,"Franche-Comté"
"Y_GE25","FR5",2006,5.9,"Ouest (FR)"
"Y_GE25","FR51",2006,5.6,"Pays de la Loire"
"Y_GE25","FR52",2006,6,"Bretagne"
"Y_GE25","FR53",2006,6.2,"Poitou-Charentes"
"Y_GE25","FR6",2006,6.4,"Sud-Ouest (FR)"
"Y_GE25","FR61",2006,6.2,"Aquitaine"
"Y_GE25","FR62",2006,7.2,"Midi-Pyrénées"
"Y_GE25","FR63",2006,4.4,"Limousin"
"Y_GE25","FR7",2006,5.8,"Centre-Est (FR)"
"Y_GE25","FR71",2006,5.8,"Rhône-Alpes"
"Y_GE25","FR72",2006,5.9,"Auvergne"
"Y_GE25","FR8",2006,9.2,"Méditerranée"
"Y_GE25","FR81",2006,9,"Languedoc-Roussillon"
"Y_GE25","FR82",2006,9.3,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2006,9.5,"Corse"
"Y_GE25","FR9",2006,23.3,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2006,23.7,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2006,20.9,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2006,26.1,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2006,23.9,"Réunion (NUTS 2010)"
"Y_GE25","HR",2006,9,"Croatia"
"Y_GE25","HR0",2006,9,"Hrvatska"
"Y_GE25","HU",2006,6.5,"Hungary"
"Y_GE25","HU1",2006,4.5,"Közép-Magyarország"
"Y_GE25","HU10",2006,4.5,"Közép-Magyarország"
"Y_GE25","HU2",2006,6,"Dunántúl"
"Y_GE25","HU21",2006,5.3,"Közép-Dunántúl"
"Y_GE25","HU22",2006,5.1,"Nyugat-Dunántúl"
"Y_GE25","HU23",2006,8.1,"Dél-Dunántúl"
"Y_GE25","HU3",2006,8.6,"Alföld és Észak"
"Y_GE25","HU31",2006,9.5,"Észak-Magyarország"
"Y_GE25","HU32",2006,9.3,"Észak-Alföld"
"Y_GE25","HU33",2006,6.9,"Dél-Alföld"
"Y_GE25","IE",2006,3.6,"Ireland"
"Y_GE25","IE0",2006,3.6,"Éire/Ireland"
"Y_GE25","IE01",2006,3.6,"Border, Midland and Western"
"Y_GE25","IE02",2006,3.6,"Southern and Eastern"
"Y_GE25","IS",2006,1.7,"Iceland"
"Y_GE25","IS0",2006,1.7,"Ísland"
"Y_GE25","IS00",2006,1.7,"Ísland"
"Y_GE25","IT",2006,5.5,"Italy"
"Y_GE25","ITC",2006,3.2,"Nord-Ovest"
"Y_GE25","ITC1",2006,3.2,"Piemonte"
"Y_GE25","ITC2",2006,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2006,4.1,"Liguria"
"Y_GE25","ITC4",2006,3,"Lombardia"
"Y_GE25","ITF",2006,9.7,"Sud"
"Y_GE25","ITF1",2006,5.5,"Abruzzo"
"Y_GE25","ITF2",2006,8.4,"Molise"
"Y_GE25","ITF3",2006,10.3,"Campania"
"Y_GE25","ITF4",2006,10.2,"Puglia"
"Y_GE25","ITF5",2006,8.7,"Basilicata"
"Y_GE25","ITF6",2006,10.7,"Calabria"
"Y_GE25","ITG",2006,10.1,"Isole"
"Y_GE25","ITG1",2006,10.6,"Sicilia"
"Y_GE25","ITG2",2006,8.8,"Sardegna"
"Y_GE25","ITH",2006,3,"Nord-Est"
"Y_GE25","ITH1",2006,2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2006,2.6,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2006,3.4,"Veneto"
"Y_GE25","ITH4",2006,2.9,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2006,2.9,"Emilia-Romagna"
"Y_GE25","ITI",2006,5.1,"Centro (IT)"
"Y_GE25","ITI1",2006,4.1,"Toscana"
"Y_GE25","ITI2",2006,4.3,"Umbria"
"Y_GE25","ITI3",2006,4,"Marche"
"Y_GE25","ITI4",2006,6.2,"Lazio"
"Y_GE25","LT",2006,5.4,"Lithuania"
"Y_GE25","LT0",2006,5.4,"Lietuva"
"Y_GE25","LT00",2006,5.4,"Lietuva"
"Y_GE25","LU",2006,3.9,"Luxembourg"
"Y_GE25","LU0",2006,3.9,"Luxembourg"
"Y_GE25","LU00",2006,3.9,"Luxembourg"
"Y_GE25","LV",2006,6.1,"Latvia"
"Y_GE25","LV0",2006,6.1,"Latvija"
"Y_GE25","LV00",2006,6.1,"Latvija"
"Y_GE25","MK",2006,32.5,"Former Yugoslav Republic of Macedonia, the"
"Y_GE25","MK0",2006,32.5,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MK00",2006,32.5,"Poranesna jugoslovenska Republika Makedonija"
"Y_GE25","MT",2006,4.8,"Malta"
"Y_GE25","MT0",2006,4.8,"Malta"
"Y_GE25","MT00",2006,4.8,"Malta"
"Y_GE25","NL",2006,3.4,"Netherlands"
"Y_GE25","NL1",2006,3.9,"Noord-Nederland"
"Y_GE25","NL11",2006,4.4,"Groningen"
"Y_GE25","NL12",2006,3.7,"Friesland (NL)"
"Y_GE25","NL13",2006,3.7,"Drenthe"
"Y_GE25","NL2",2006,3.3,"Oost-Nederland"
"Y_GE25","NL21",2006,3.6,"Overijssel"
"Y_GE25","NL22",2006,2.9,"Gelderland"
"Y_GE25","NL23",2006,4.2,"Flevoland"
"Y_GE25","NL3",2006,3.4,"West-Nederland"
"Y_GE25","NL31",2006,2.8,"Utrecht"
"Y_GE25","NL32",2006,3.4,"Noord-Holland"
"Y_GE25","NL33",2006,3.7,"Zuid-Holland"
"Y_GE25","NL34",2006,2.4,"Zeeland"
"Y_GE25","NL4",2006,3.3,"Zuid-Nederland"
"Y_GE25","NL41",2006,3,"Noord-Brabant"
"Y_GE25","NL42",2006,3.9,"Limburg (NL)"
"Y_GE25","NO",2006,2.6,"Norway"
"Y_GE25","NO0",2006,2.6,"Norge"
"Y_GE25","NO01",2006,2.9,"Oslo og Akershus"
"Y_GE25","NO02",2006,2.1,"Hedmark og Oppland"
"Y_GE25","NO03",2006,3,"Sør-Østlandet"
"Y_GE25","NO04",2006,2.2,"Agder og Rogaland"
"Y_GE25","NO05",2006,2,"Vestlandet"
"Y_GE25","NO06",2006,2.6,"Trøndelag"
"Y_GE25","NO07",2006,2.7,"Nord-Norge"
"Y_GE25","PL",2006,11.7,"Poland"
"Y_GE25","PL1",2006,11,"Region Centralny"
"Y_GE25","PL11",2006,12.1,"Lódzkie"
"Y_GE25","PL12",2006,10.4,"Mazowieckie"
"Y_GE25","PL2",2006,11.2,"Region Poludniowy"
"Y_GE25","PL21",2006,10.1,"Malopolskie"
"Y_GE25","PL22",2006,12.1,"Slaskie"
"Y_GE25","PL3",2006,10.8,"Region Wschodni"
"Y_GE25","PL31",2006,10.1,"Lubelskie"
"Y_GE25","PL32",2006,11,"Podkarpackie"
"Y_GE25","PL33",2006,12.6,"Swietokrzyskie"
"Y_GE25","PL34",2006,9.4,"Podlaskie"
"Y_GE25","PL4",2006,12,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2006,10.4,"Wielkopolskie"
"Y_GE25","PL42",2006,15.5,"Zachodniopomorskie"
"Y_GE25","PL43",2006,12.2,"Lubuskie"
"Y_GE25","PL5",2006,14.4,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2006,15.4,"Dolnoslaskie"
"Y_GE25","PL52",2006,11.3,"Opolskie"
"Y_GE25","PL6",2006,13.2,"Region Pólnocny"
"Y_GE25","PL61",2006,13.9,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2006,14,"Warminsko-Mazurskie"
"Y_GE25","PL63",2006,11.8,"Pomorskie"
"Y_GE25","PT",2006,6.7,"Portugal"
"Y_GE25","PT1",2006,6.9,"Continente"
"Y_GE25","PT11",2006,7.9,"Norte"
"Y_GE25","PT15",2006,4.7,"Algarve"
"Y_GE25","PT16",2006,4.8,"Centro (PT)"
"Y_GE25","PT17",2006,7.5,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2006,7.8,"Alentejo"
"Y_GE25","PT2",2006,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2006,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2006,4.6,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2006,4.6,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2006,5.7,"Romania"
"Y_GE25","RO1",2006,5.9,"Macroregiunea unu"
"Y_GE25","RO11",2006,4.6,"Nord-Vest"
"Y_GE25","RO12",2006,7.4,"Centru"
"Y_GE25","RO2",2006,5.6,"Macroregiunea doi"
"Y_GE25","RO21",2006,4.5,"Nord-Est"
"Y_GE25","RO22",2006,7.1,"Sud-Est"
"Y_GE25","RO3",2006,5.8,"Macroregiunea trei"
"Y_GE25","RO31",2006,7.1,"Sud - Muntenia"
"Y_GE25","RO32",2006,3.9,"Bucuresti - Ilfov"
"Y_GE25","RO4",2006,5.6,"Macroregiunea patru"
"Y_GE25","RO41",2006,5.6,"Sud-Vest Oltenia"
"Y_GE25","RO42",2006,5.5,"Vest"
"Y_GE25","SE",2006,5,"Sweden"
"Y_GE25","SE1",2006,4.8,"Östra Sverige"
"Y_GE25","SE11",2006,4.6,"Stockholm"
"Y_GE25","SE12",2006,5.2,"Östra Mellansverige"
"Y_GE25","SE2",2006,4.9,"Södra Sverige"
"Y_GE25","SE21",2006,4.1,"Småland med öarna"
"Y_GE25","SE22",2006,5.8,"Sydsverige"
"Y_GE25","SE23",2006,4.7,"Västsverige"
"Y_GE25","SE3",2006,5.8,"Norra Sverige"
"Y_GE25","SE31",2006,5.7,"Norra Mellansverige"
"Y_GE25","SE32",2006,5.7,"Mellersta Norrland"
"Y_GE25","SE33",2006,6.1,"Övre Norrland"
"Y_GE25","SI",2006,5,"Slovenia"
"Y_GE25","SI0",2006,5,"Slovenija"
"Y_GE25","SI01",2006,5.9,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2006,4,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2006,11.7,"Slovakia"
"Y_GE25","SK0",2006,11.7,"Slovensko"
"Y_GE25","SK01",2006,4.2,"Bratislavský kraj"
"Y_GE25","SK02",2006,8.4,"Západné Slovensko"
"Y_GE25","SK03",2006,14.7,"Stredné Slovensko"
"Y_GE25","SK04",2006,16.7,"Východné Slovensko"
"Y_GE25","TR",2006,6.9,"Turkey"
"Y_GE25","TR1",2006,9,"Istanbul"
"Y_GE25","TR10",2006,9,"Istanbul"
"Y_GE25","TR2",2006,4.2,"Bati Marmara"
"Y_GE25","TR21",2006,5,"Tekirdag, Edirne, Kirklareli"
"Y_GE25","TR22",2006,3.5,"Balikesir, Çanakkale"
"Y_GE25","TR3",2006,5.9,"Ege"
"Y_GE25","TR31",2006,8.4,"Izmir"
"Y_GE25","TR32",2006,4.1,"Aydin, Denizli, Mugla"
"Y_GE25","TR33",2006,4.7,"Manisa, Afyonkarahisar, Kütahya, Usak"
"Y_GE25","TR4",2006,6.7,"Dogu Marmara"
"Y_GE25","TR41",2006,5.4,"Bursa, Eskisehir, Bilecik"
"Y_GE25","TR42",2006,8.2,"Kocaeli, Sakarya, Düzce, Bolu, Yalova"
"Y_GE25","TR5",2006,8.3,"Bati Anadolu"
"Y_GE25","TR51",2006,8.9,"Ankara"
"Y_GE25","TR52",2006,6.8,"Konya, Karaman"
"Y_GE25","TR6",2006,8.7,"Akdeniz"
"Y_GE25","TR61",2006,5.2,"Antalya, Isparta, Burdur"
"Y_GE25","TR62",2006,11.8,"Adana, Mersin"
"Y_GE25","TR63",2006,8.4,"Hatay, Kahramanmaras, Osmaniye"
"Y_GE25","TR7",2006,6.6,"Orta Anadolu"
"Y_GE25","TR71",2006,6.7,"Kirikkale, Aksaray, Nigde, Nevsehir, Kirsehir"
"Y_GE25","TR72",2006,6.6,"Kayseri, Sivas, Yozgat"
"Y_GE25","TR8",2006,3.8,"Bati Karadeniz"
"Y_GE25","TR81",2006,3.1,"Zonguldak, Karabük, Bartin"
"Y_GE25","TR82",2006,2.6,"Kastamonu, Çankiri, Sinop"
"Y_GE25","TR83",2006,4.5,"Samsun, Tokat, Çorum, Amasya"
"Y_GE25","TR9",2006,2.7,"Dogu Karadeniz"
"Y_GE25","TR90",2006,2.7,"Trabzon, Ordu, Giresun, Rize, Artvin, Gümüshane"
"Y_GE25","TRA",2006,2.6,"Kuzeydogu Anadolu"
"Y_GE25","TRA1",2006,3.1,"Erzurum, Erzincan, Bayburt"
"Y_GE25","TRA2",2006,2.1,"Agri, Kars, Igdir, Ardahan"
"Y_GE25","TRB",2006,6.7,"Ortadogu Anadolu"
"Y_GE25","TRB1",2006,7.5,"Malatya, Elazig, Bingöl, Tunceli"
"Y_GE25","TRB2",2006,5.6,"Van, Mus, Bitlis, Hakkari"
"Y_GE25","TRC",2006,10.3,"Güneydogu Anadolu"
"Y_GE25","TRC1",2006,11.2,"Gaziantep, Adiyaman, Kilis"
"Y_GE25","TRC2",2006,8.8,"Sanliurfa, Diyarbakir"
"Y_GE25","TRC3",2006,11.1,"Mardin, Batman, Sirnak, Siirt"
"Y_GE25","UK",2006,3.8,"United Kingdom"
"Y_GE25","UKC",2006,4.6,"North East (UK)"
"Y_GE25","UKC1",2006,3.7,"Tees Valley and Durham"
"Y_GE25","UKC2",2006,5.3,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2006,3.4,"North West (UK)"
"Y_GE25","UKD1",2006,2.9,"Cumbria"
"Y_GE25","UKD3",2006,3.8,"Greater Manchester"
"Y_GE25","UKD4",2006,2.9,"Lancashire"
"Y_GE25","UKD6",2006,2.5,"Cheshire"
"Y_GE25","UKD7",2006,4.2,"Merseyside"
"Y_GE25","UKE",2006,3.9,"Yorkshire and The Humber"
"Y_GE25","UKE1",2006,4.1,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2006,2.6,"North Yorkshire"
"Y_GE25","UKE3",2006,4.9,"South Yorkshire"
"Y_GE25","UKE4",2006,3.6,"West Yorkshire"
"Y_GE25","UKF",2006,3.4,"East Midlands (UK)"
"Y_GE25","UKF1",2006,3.6,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2006,3.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2006,3.2,"Lincolnshire"
"Y_GE25","UKG",2006,3.9,"West Midlands (UK)"
"Y_GE25","UKG1",2006,2.5,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2006,2.7,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2006,5.6,"West Midlands"
"Y_GE25","UKH",2006,3.5,"East of England"
"Y_GE25","UKH1",2006,3.4,"East Anglia"
"Y_GE25","UKH2",2006,3.5,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2006,3.4,"Essex"
"Y_GE25","UKI",2006,5.9,"London"
"Y_GE25","UKI1",2006,7.1,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2006,5.1,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2006,3.2,"South East (UK)"
"Y_GE25","UKJ1",2006,2.6,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2006,3.1,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2006,3.4,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2006,3.8,"Kent"
"Y_GE25","UKK",2006,2.6,"South West (UK)"
"Y_GE25","UKK1",2006,2.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2006,3,"Dorset and Somerset"
"Y_GE25","UKK3",2006,2.9,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2006,2.7,"Devon"
"Y_GE25","UKL",2006,3.5,"Wales"
"Y_GE25","UKL1",2006,3.5,"West Wales and The Valleys"
"Y_GE25","UKL2",2006,3.6,"East Wales"
"Y_GE25","UKM",2006,3.6,"Scotland"
"Y_GE25","UKM2",2006,3.4,"Eastern Scotland"
"Y_GE25","UKM3",2006,4.5,"South Western Scotland"
"Y_GE25","UKM5",2006,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2006,2.4,"Highlands and Islands"
"Y_GE25","UKN",2006,3.3,"Northern Ireland (UK)"
"Y_GE25","UKN0",2006,3.3,"Northern Ireland (UK)"
"Y15-24","AT",2005,11,"Austria"
"Y15-24","AT1",2005,15,"Ostösterreich"
"Y15-24","AT11",2005,NA,"Burgenland (AT)"
"Y15-24","AT12",2005,9.7,"Niederösterreich"
"Y15-24","AT13",2005,21.2,"Wien"
"Y15-24","AT2",2005,9.3,"Südösterreich"
"Y15-24","AT21",2005,10.9,"Kärnten"
"Y15-24","AT22",2005,8.6,"Steiermark"
"Y15-24","AT3",2005,8.2,"Westösterreich"
"Y15-24","AT31",2005,7.4,"Oberösterreich"
"Y15-24","AT32",2005,7.8,"Salzburg"
"Y15-24","AT33",2005,8.9,"Tirol"
"Y15-24","AT34",2005,10.6,"Vorarlberg"
"Y15-24","BE",2005,21.5,"Belgium"
"Y15-24","BE1",2005,35.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2005,35.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2005,14.2,"Vlaams Gewest"
"Y15-24","BE21",2005,11.8,"Prov. Antwerpen"
"Y15-24","BE22",2005,16.1,"Prov. Limburg (BE)"
"Y15-24","BE23",2005,16.6,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2005,16.1,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2005,11.9,"Prov. West-Vlaanderen"
"Y15-24","BE3",2005,31.8,"Région wallonne"
"Y15-24","BE31",2005,28.8,"Prov. Brabant Wallon"
"Y15-24","BE32",2005,36.6,"Prov. Hainaut"
"Y15-24","BE33",2005,28,"Prov. Liège"
"Y15-24","BE34",2005,23.7,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2005,32.6,"Prov. Namur"
"Y15-24","BG",2005,22.3,"Bulgaria"
"Y15-24","BG3",2005,24.6,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2005,30.8,"Severozapaden"
"Y15-24","BG32",2005,25.6,"Severen tsentralen"
"Y15-24","BG33",2005,25.1,"Severoiztochen"
"Y15-24","BG34",2005,18.9,"Yugoiztochen"
"Y15-24","BG4",2005,20.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2005,14.7,"Yugozapaden"
"Y15-24","BG42",2005,28.8,"Yuzhen tsentralen"
"Y15-24","CH",2005,8.8,"Switzerland"
"Y15-24","CH0",2005,8.8,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2005,13.8,"Région lémanique"
"Y15-24","CH02",2005,8.1,"Espace Mittelland"
"Y15-24","CH03",2005,7.5,"Nordwestschweiz"
"Y15-24","CH04",2005,6.8,"Zürich"
"Y15-24","CH05",2005,8.7,"Ostschweiz"
"Y15-24","CH06",2005,5.5,"Zentralschweiz"
"Y15-24","CH07",2005,15.8,"Ticino"
"Y15-24","CY",2005,13.9,"Cyprus"
"Y15-24","CY0",2005,13.9,"Kypros"
"Y15-24","CY00",2005,13.9,"Kypros"
"Y15-24","CZ",2005,19.2,"Czech Republic"
"Y15-24","CZ0",2005,19.2,"Ceská republika"
"Y15-24","CZ01",2005,9.2,"Praha"
"Y15-24","CZ02",2005,11.1,"Strední Cechy"
"Y15-24","CZ03",2005,12.4,"Jihozápad"
"Y15-24","CZ04",2005,27.8,"Severozápad"
"Y15-24","CZ05",2005,14.8,"Severovýchod"
"Y15-24","CZ06",2005,19.9,"Jihovýchod"
"Y15-24","CZ07",2005,22.4,"Strední Morava"
"Y15-24","CZ08",2005,32.2,"Moravskoslezsko"
"Y15-24","DE",2005,15.5,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2005,11.1,"Baden-Württemberg"
"Y15-24","DE11",2005,10.8,"Stuttgart"
"Y15-24","DE12",2005,11.9,"Karlsruhe"
"Y15-24","DE13",2005,10.6,"Freiburg"
"Y15-24","DE14",2005,11.2,"Tübingen"
"Y15-24","DE2",2005,11.6,"Bayern"
"Y15-24","DE21",2005,10.4,"Oberbayern"
"Y15-24","DE22",2005,9.2,"Niederbayern"
"Y15-24","DE23",2005,10.2,"Oberpfalz"
"Y15-24","DE24",2005,16.4,"Oberfranken"
"Y15-24","DE25",2005,13.1,"Mittelfranken"
"Y15-24","DE26",2005,16,"Unterfranken"
"Y15-24","DE27",2005,9.4,"Schwaben"
"Y15-24","DE3",2005,23.9,"Berlin"
"Y15-24","DE30",2005,23.9,"Berlin"
"Y15-24","DE4",2005,22.5,"Brandenburg"
"Y15-24","DE40",2005,22.5,"Brandenburg"
"Y15-24","DE5",2005,19.3,"Bremen"
"Y15-24","DE50",2005,19.3,"Bremen"
"Y15-24","DE6",2005,14.7,"Hamburg"
"Y15-24","DE60",2005,14.7,"Hamburg"
"Y15-24","DE7",2005,13,"Hessen"
"Y15-24","DE71",2005,12.1,"Darmstadt"
"Y15-24","DE72",2005,16.1,"Gießen"
"Y15-24","DE73",2005,12.4,"Kassel"
"Y15-24","DE8",2005,20.9,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2005,20.9,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2005,16.2,"Niedersachsen"
"Y15-24","DE91",2005,19.1,"Braunschweig"
"Y15-24","DE92",2005,16.8,"Hannover"
"Y15-24","DE93",2005,15.9,"Lüneburg"
"Y15-24","DE94",2005,14.2,"Weser-Ems"
"Y15-24","DEA",2005,15.6,"Nordrhein-Westfalen"
"Y15-24","DEA1",2005,15.4,"Düsseldorf"
"Y15-24","DEA2",2005,14.7,"Köln"
"Y15-24","DEA3",2005,15.1,"Münster"
"Y15-24","DEA4",2005,15.2,"Detmold"
"Y15-24","DEA5",2005,17.5,"Arnsberg"
"Y15-24","DEB",2005,13.8,"Rheinland-Pfalz"
"Y15-24","DEB1",2005,13.9,"Koblenz"
"Y15-24","DEB2",2005,NA,"Trier"
"Y15-24","DEB3",2005,14.4,"Rheinhessen-Pfalz"
"Y15-24","DEC",2005,17.8,"Saarland"
"Y15-24","DEC0",2005,17.8,"Saarland"
"Y15-24","DED",2005,20.4,"Sachsen"
"Y15-24","DED2",2005,20.7,"Dresden"
"Y15-24","DED4",2005,17.1,"Chemnitz"
"Y15-24","DED5",2005,24.7,"Leipzig"
"Y15-24","DEE",2005,23.4,"Sachsen-Anhalt"
"Y15-24","DEE0",2005,23.4,"Sachsen-Anhalt"
"Y15-24","DEF",2005,15.5,"Schleswig-Holstein"
"Y15-24","DEF0",2005,15.5,"Schleswig-Holstein"
"Y15-24","DEG",2005,19.3,"Thüringen"
"Y15-24","DEG0",2005,19.3,"Thüringen"
"Y15-24","DK",2005,8.6,"Denmark"
"Y15-24","DK0",2005,8.6,"Danmark"
"Y15-24","EA17",2005,18.1,"Euro area (17 countries)"
"Y15-24","EA18",2005,18,"Euro area (18 countries)"
"Y15-24","EA19",2005,18,"Euro area (19 countries)"
"Y15-24","EE",2005,15.1,"Estonia"
"Y15-24","EE0",2005,15.1,"Eesti"
"Y15-24","EE00",2005,15.1,"Eesti"
"Y15-24","EL",2005,25.8,"Greece"
"Y15-24","EL1",2005,28.7,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2005,31.3,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2005,28.7,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2005,44.4,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2005,20,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2005,29.2,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2005,36.3,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2005,23.7,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2005,25,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2005,31.4,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2005,30.9,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2005,23,"Attiki"
"Y15-24","EL30",2005,23,"Attiki"
"Y15-24","EL4",2005,21.4,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2005,37.3,"Voreio Aigaio"
"Y15-24","EL42",2005,18.3,"Notio Aigaio"
"Y15-24","EL43",2005,17.8,"Kriti"
"Y15-24","ES",2005,19.6,"Spain"
"Y15-24","ES1",2005,21,"Noroeste (ES)"
"Y15-24","ES11",2005,20.8,"Galicia"
"Y15-24","ES12",2005,23.7,"Principado de Asturias"
"Y15-24","ES13",2005,17.9,"Cantabria"
"Y15-24","ES2",2005,16,"Noreste (ES)"
"Y15-24","ES21",2005,18.9,"País Vasco"
"Y15-24","ES22",2005,14.7,"Comunidad Foral de Navarra"
"Y15-24","ES23",2005,14.4,"La Rioja"
"Y15-24","ES24",2005,13,"Aragón"
"Y15-24","ES3",2005,16.7,"Comunidad de Madrid"
"Y15-24","ES30",2005,16.7,"Comunidad de Madrid"
"Y15-24","ES4",2005,20.9,"Centro (ES)"
"Y15-24","ES41",2005,19.4,"Castilla y León"
"Y15-24","ES42",2005,18.2,"Castilla-la Mancha"
"Y15-24","ES43",2005,28.6,"Extremadura"
"Y15-24","ES5",2005,17.4,"Este (ES)"
"Y15-24","ES51",2005,15.8,"Cataluña"
"Y15-24","ES52",2005,19.6,"Comunidad Valenciana"
"Y15-24","ES53",2005,18.2,"Illes Balears"
"Y15-24","ES6",2005,23.4,"Sur (ES)"
"Y15-24","ES61",2005,24.6,"Andalucía"
"Y15-24","ES62",2005,15.4,"Región de Murcia"
"Y15-24","ES63",2005,44.5,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2005,38.1,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2005,24.4,"Canarias (ES)"
"Y15-24","ES70",2005,24.4,"Canarias (ES)"
"Y15-24","EU15",2005,16.7,"European Union (15 countries)"
"Y15-24","EU27",2005,18.7,"European Union (27 countries)"
"Y15-24","EU28",2005,18.8,"European Union (28 countries)"
"Y15-24","FI",2005,20.1,"Finland"
"Y15-24","FI1",2005,20.1,"Manner-Suomi"
"Y15-24","FI19",2005,20.8,"Länsi-Suomi"
"Y15-24","FI1B",2005,15.5,"Helsinki-Uusimaa"
"Y15-24","FI1C",2005,19.2,"Etelä-Suomi"
"Y15-24","FI1D",2005,26,"Pohjois- ja Itä-Suomi"
"Y15-24","FI2",2005,NA,"Åland"
"Y15-24","FI20",2005,NA,"Åland"
"Y15-24","FR",2005,21.1,"France"
"Y15-24","FR1",2005,18.6,"Île de France"
"Y15-24","FR10",2005,18.6,"Île de France"
"Y15-24","FR2",2005,21.8,"Bassin Parisien"
"Y15-24","FR21",2005,21.9,"Champagne-Ardenne"
"Y15-24","FR22",2005,29.7,"Picardie"
"Y15-24","FR23",2005,18.2,"Haute-Normandie"
"Y15-24","FR24",2005,20.9,"Centre (FR)"
"Y15-24","FR25",2005,21.6,"Basse-Normandie"
"Y15-24","FR26",2005,19.4,"Bourgogne"
"Y15-24","FR3",2005,29.4,"Nord - Pas-de-Calais"
"Y15-24","FR30",2005,29.4,"Nord - Pas-de-Calais"
"Y15-24","FR4",2005,20.5,"Est (FR)"
"Y15-24","FR41",2005,23.9,"Lorraine"
"Y15-24","FR42",2005,18.2,"Alsace"
"Y15-24","FR43",2005,17,"Franche-Comté"
"Y15-24","FR5",2005,18.5,"Ouest (FR)"
"Y15-24","FR51",2005,19.4,"Pays de la Loire"
"Y15-24","FR52",2005,15.9,"Bretagne"
"Y15-24","FR53",2005,21.1,"Poitou-Charentes"
"Y15-24","FR6",2005,16.1,"Sud-Ouest (FR)"
"Y15-24","FR61",2005,17.2,"Aquitaine"
"Y15-24","FR62",2005,14.4,"Midi-Pyrénées"
"Y15-24","FR63",2005,NA,"Limousin"
"Y15-24","FR7",2005,16.8,"Centre-Est (FR)"
"Y15-24","FR71",2005,17.1,"Rhône-Alpes"
"Y15-24","FR72",2005,15.9,"Auvergne"
"Y15-24","FR8",2005,23.6,"Méditerranée"
"Y15-24","FR81",2005,25.5,"Languedoc-Roussillon"
"Y15-24","FR82",2005,22.5,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2005,NA,"Corse"
"Y15-24","FR9",2005,51.9,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2005,59.1,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2005,42.7,"Martinique (NUTS 2010)"
"Y15-24","FR93",2005,52.5,"Guyane (NUTS 2010)"
"Y15-24","FR94",2005,52.2,"Réunion (NUTS 2010)"
"Y15-24","HR",2005,32.3,"Croatia"
"Y15-24","HR0",2005,32.3,"Hrvatska"
"Y15-24","HU",2005,19.4,"Hungary"
"Y15-24","HU1",2005,14.4,"Közép-Magyarország"
"Y15-24","HU10",2005,14.4,"Közép-Magyarország"
"Y15-24","HU2",2005,16.8,"Dunántúl"
"Y15-24","HU21",2005,13.9,"Közép-Dunántúl"
"Y15-24","HU22",2005,13.5,"Nyugat-Dunántúl"
"Y15-24","HU23",2005,24.9,"Dél-Dunántúl"
"Y15-24","HU3",2005,24.7,"Alföld és Észak"
"Y15-24","HU31",2005,28.5,"Észak-Magyarország"
"Y15-24","HU32",2005,24.8,"Észak-Alföld"
"Y15-24","HU33",2005,21,"Dél-Alföld"
"Y15-24","IE",2005,8.6,"Ireland"
"Y15-24","IE0",2005,8.6,"Éire/Ireland"
"Y15-24","IE01",2005,8.7,"Border, Midland and Western"
"Y15-24","IE02",2005,8.5,"Southern and Eastern"
"Y15-24","IS",2005,7.4,"Iceland"
"Y15-24","IS0",2005,7.4,"Ísland"
"Y15-24","IS00",2005,7.4,"Ísland"
"Y15-24","IT",2005,24.1,"Italy"
"Y15-24","ITC",2005,14.8,"Nord-Ovest"
"Y15-24","ITC1",2005,17,"Piemonte"
"Y15-24","ITC2",2005,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2005,19.9,"Liguria"
"Y15-24","ITC4",2005,13.2,"Lombardia"
"Y15-24","ITF",2005,37.4,"Sud"
"Y15-24","ITF1",2005,23.1,"Abruzzo"
"Y15-24","ITF2",2005,31.3,"Molise"
"Y15-24","ITF3",2005,39,"Campania"
"Y15-24","ITF4",2005,35.7,"Puglia"
"Y15-24","ITF5",2005,36.5,"Basilicata"
"Y15-24","ITF6",2005,46.1,"Calabria"
"Y15-24","ITG",2005,41.5,"Isole"
"Y15-24","ITG1",2005,44.8,"Sicilia"
"Y15-24","ITG2",2005,32.6,"Sardegna"
"Y15-24","ITH",2005,11.5,"Nord-Est"
"Y15-24","ITH1",2005,7.2,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2005,10.4,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2005,12.6,"Veneto"
"Y15-24","ITH4",2005,10.6,"Friuli-Venezia Giulia"
"Y15-24","ITH5",2005,11.3,"Emilia-Romagna"
"Y15-24","ITI",2005,21.2,"Centro (IT)"
"Y15-24","ITI1",2005,16.9,"Toscana"
"Y15-24","ITI2",2005,18.2,"Umbria"
"Y15-24","ITI3",2005,15.2,"Marche"
"Y15-24","ITI4",2005,26.7,"Lazio"
"Y15-24","LT",2005,15.8,"Lithuania"
"Y15-24","LT0",2005,15.8,"Lietuva"
"Y15-24","LT00",2005,15.8,"Lietuva"
"Y15-24","LU",2005,13.7,"Luxembourg"
"Y15-24","LU0",2005,13.7,"Luxembourg"
"Y15-24","LU00",2005,13.7,"Luxembourg"
"Y15-24","LV",2005,15.1,"Latvia"
"Y15-24","LV0",2005,15.1,"Latvija"
"Y15-24","LV00",2005,15.1,"Latvija"
"Y15-24","MT",2005,16.1,"Malta"
"Y15-24","MT0",2005,16.1,"Malta"
"Y15-24","MT00",2005,16.1,"Malta"
"Y15-24","NL",2005,8.2,"Netherlands"
"Y15-24","NL1",2005,9.8,"Noord-Nederland"
"Y15-24","NL11",2005,9.7,"Groningen"
"Y15-24","NL12",2005,9.6,"Friesland (NL)"
"Y15-24","NL13",2005,10.3,"Drenthe"
"Y15-24","NL2",2005,8.2,"Oost-Nederland"
"Y15-24","NL21",2005,7.9,"Overijssel"
"Y15-24","NL22",2005,7.7,"Gelderland"
"Y15-24","NL23",2005,11.2,"Flevoland"
"Y15-24","NL3",2005,8.4,"West-Nederland"
"Y15-24","NL31",2005,6.8,"Utrecht"
"Y15-24","NL32",2005,8.1,"Noord-Holland"
"Y15-24","NL33",2005,9.4,"Zuid-Holland"
"Y15-24","NL34",2005,6.2,"Zeeland"
"Y15-24","NL4",2005,7,"Zuid-Nederland"
"Y15-24","NL41",2005,6.5,"Noord-Brabant"
"Y15-24","NL42",2005,8.3,"Limburg (NL)"
"Y15-24","NO",2005,11.5,"Norway"
"Y15-24","NO0",2005,11.5,"Norge"
"Y15-24","NO01",2005,10.7,"Oslo og Akershus"
"Y15-24","NO02",2005,12,"Hedmark og Oppland"
"Y15-24","NO03",2005,12.3,"Sør-Østlandet"
"Y15-24","NO04",2005,11.1,"Agder og Rogaland"
"Y15-24","NO05",2005,10.5,"Vestlandet"
"Y15-24","NO06",2005,10.2,"Trøndelag"
"Y15-24","NO07",2005,14.6,"Nord-Norge"
"Y15-24","PL",2005,36.9,"Poland"
"Y15-24","PL1",2005,32.3,"Region Centralny"
"Y15-24","PL11",2005,33.1,"Lódzkie"
"Y15-24","PL12",2005,31.9,"Mazowieckie"
"Y15-24","PL2",2005,38,"Region Poludniowy"
"Y15-24","PL21",2005,36.7,"Malopolskie"
"Y15-24","PL22",2005,38.8,"Slaskie"
"Y15-24","PL3",2005,36.5,"Region Wschodni"
"Y15-24","PL31",2005,30.3,"Lubelskie"
"Y15-24","PL32",2005,43.3,"Podkarpackie"
"Y15-24","PL33",2005,43.6,"Swietokrzyskie"
"Y15-24","PL34",2005,30.6,"Podlaskie"
"Y15-24","PL4",2005,36.5,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2005,34.9,"Wielkopolskie"
"Y15-24","PL42",2005,41.7,"Zachodniopomorskie"
"Y15-24","PL43",2005,35.3,"Lubuskie"
"Y15-24","PL5",2005,42.8,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2005,45,"Dolnoslaskie"
"Y15-24","PL52",2005,36.1,"Opolskie"
"Y15-24","PL6",2005,38.2,"Region Pólnocny"
"Y15-24","PL61",2005,39.1,"Kujawsko-Pomorskie"
"Y15-24","PL62",2005,39.9,"Warminsko-Mazurskie"
"Y15-24","PL63",2005,36.3,"Pomorskie"
"Y15-24","PT",2005,16.2,"Portugal"
"Y15-24","PT1",2005,16.6,"Continente"
"Y15-24","PT11",2005,16.1,"Norte"
"Y15-24","PT15",2005,NA,"Algarve"
"Y15-24","PT16",2005,14.8,"Centro (PT)"
"Y15-24","PT17",2005,18.3,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2005,20.7,"Alentejo"
"Y15-24","PT2",2005,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2005,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2005,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2005,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2005,20.2,"Romania"
"Y15-24","RO1",2005,19.3,"Macroregiunea unu"
"Y15-24","RO11",2005,18.8,"Nord-Vest"
"Y15-24","RO12",2005,19.9,"Centru"
"Y15-24","RO2",2005,18.5,"Macroregiunea doi"
"Y15-24","RO21",2005,17.1,"Nord-Est"
"Y15-24","RO22",2005,20.6,"Sud-Est"
"Y15-24","RO3",2005,24.4,"Macroregiunea trei"
"Y15-24","RO31",2005,25,"Sud - Muntenia"
"Y15-24","RO32",2005,23.4,"Bucuresti - Ilfov"
"Y15-24","RO4",2005,18.8,"Macroregiunea patru"
"Y15-24","RO41",2005,19.1,"Sud-Vest Oltenia"
"Y15-24","RO42",2005,18.5,"Vest"
"Y15-24","SE",2005,22.8,"Sweden"
"Y15-24","SE1",2005,22,"Östra Sverige"
"Y15-24","SE11",2005,21.5,"Stockholm"
"Y15-24","SE12",2005,22.7,"Östra Mellansverige"
"Y15-24","SE2",2005,22.4,"Södra Sverige"
"Y15-24","SE21",2005,18.9,"Småland med öarna"
"Y15-24","SE22",2005,22.3,"Sydsverige"
"Y15-24","SE23",2005,24.1,"Västsverige"
"Y15-24","SE3",2005,25.4,"Norra Sverige"
"Y15-24","SE31",2005,26,"Norra Mellansverige"
"Y15-24","SE32",2005,26.4,"Mellersta Norrland"
"Y15-24","SE33",2005,24.1,"Övre Norrland"
"Y15-24","SI",2005,15.9,"Slovenia"
"Y15-24","SI0",2005,15.9,"Slovenija"
"Y15-24","SI01",2005,18.6,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2005,12.7,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2005,30.1,"Slovakia"
"Y15-24","SK0",2005,30.1,"Slovensko"
"Y15-24","SK01",2005,9.8,"Bratislavský kraj"
"Y15-24","SK02",2005,22.5,"Západné Slovensko"
"Y15-24","SK03",2005,34.7,"Stredné Slovensko"
"Y15-24","SK04",2005,41.4,"Východné Slovensko"
"Y15-24","UK",2005,12.7,"United Kingdom"
"Y15-24","UKC",2005,15.7,"North East (UK)"
"Y15-24","UKC1",2005,15.3,"Tees Valley and Durham"
"Y15-24","UKC2",2005,16,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2005,12.4,"North West (UK)"
"Y15-24","UKD1",2005,12.3,"Cumbria"
"Y15-24","UKD3",2005,12.5,"Greater Manchester"
"Y15-24","UKD4",2005,12.4,"Lancashire"
"Y15-24","UKD6",2005,8.1,"Cheshire"
"Y15-24","UKD7",2005,14.2,"Merseyside"
"Y15-24","UKE",2005,13.1,"Yorkshire and The Humber"
"Y15-24","UKE1",2005,13.9,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2005,8.3,"North Yorkshire"
"Y15-24","UKE3",2005,15.1,"South Yorkshire"
"Y15-24","UKE4",2005,13.1,"West Yorkshire"
"Y15-24","UKF",2005,11.3,"East Midlands (UK)"
"Y15-24","UKF1",2005,10.7,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2005,12.9,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2005,9.5,"Lincolnshire"
"Y15-24","UKG",2005,12.3,"West Midlands (UK)"
"Y15-24","UKG1",2005,7.8,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2005,9.2,"Shropshire and Staffordshire"
"Y15-24","UKG3",2005,15.9,"West Midlands"
"Y15-24","UKH",2005,10.7,"East of England"
"Y15-24","UKH1",2005,10.6,"East Anglia"
"Y15-24","UKH2",2005,10.5,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2005,11.1,"Essex"
"Y15-24","UKI",2005,19.7,"London"
"Y15-24","UKI1",2005,21.6,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2005,18.6,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2005,10.5,"South East (UK)"
"Y15-24","UKJ1",2005,10.7,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2005,9.3,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2005,11.4,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2005,10.8,"Kent"
"Y15-24","UKK",2005,10.1,"South West (UK)"
"Y15-24","UKK1",2005,10.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2005,7.4,"Dorset and Somerset"
"Y15-24","UKK3",2005,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2005,11.6,"Devon"
"Y15-24","UKL",2005,12.8,"Wales"
"Y15-24","UKL1",2005,14.8,"West Wales and The Valleys"
"Y15-24","UKL2",2005,9.6,"East Wales"
"Y15-24","UKM",2005,13,"Scotland"
"Y15-24","UKM2",2005,12.7,"Eastern Scotland"
"Y15-24","UKM3",2005,13.9,"South Western Scotland"
"Y15-24","UKM5",2005,12.4,"North Eastern Scotland"
"Y15-24","UKM6",2005,NA,"Highlands and Islands"
"Y15-24","UKN",2005,11.1,"Northern Ireland (UK)"
"Y15-24","UKN0",2005,11.1,"Northern Ireland (UK)"
"Y20-64","AT",2005,5.2,"Austria"
"Y20-64","AT1",2005,6.7,"Ostösterreich"
"Y20-64","AT11",2005,5.3,"Burgenland (AT)"
"Y20-64","AT12",2005,4.2,"Niederösterreich"
"Y20-64","AT13",2005,9.3,"Wien"
"Y20-64","AT2",2005,4.4,"Südösterreich"
"Y20-64","AT21",2005,4.9,"Kärnten"
"Y20-64","AT22",2005,4.2,"Steiermark"
"Y20-64","AT3",2005,3.9,"Westösterreich"
"Y20-64","AT31",2005,4.1,"Oberösterreich"
"Y20-64","AT32",2005,3.2,"Salzburg"
"Y20-64","AT33",2005,3.4,"Tirol"
"Y20-64","AT34",2005,5.2,"Vorarlberg"
"Y20-64","BE",2005,8.2,"Belgium"
"Y20-64","BE1",2005,16.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2005,16.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2005,5.3,"Vlaams Gewest"
"Y20-64","BE21",2005,6.1,"Prov. Antwerpen"
"Y20-64","BE22",2005,6.7,"Prov. Limburg (BE)"
"Y20-64","BE23",2005,4.7,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2005,4.2,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2005,4.6,"Prov. West-Vlaanderen"
"Y20-64","BE3",2005,11.4,"Région wallonne"
"Y20-64","BE31",2005,8.8,"Prov. Brabant Wallon"
"Y20-64","BE32",2005,13.4,"Prov. Hainaut"
"Y20-64","BE33",2005,11.8,"Prov. Liège"
"Y20-64","BE34",2005,7.3,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2005,10,"Prov. Namur"
"Y20-64","BG",2005,9.8,"Bulgaria"
"Y20-64","BG3",2005,10.9,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2005,12.1,"Severozapaden"
"Y20-64","BG32",2005,12.3,"Severen tsentralen"
"Y20-64","BG33",2005,11.7,"Severoiztochen"
"Y20-64","BG34",2005,7.9,"Yugoiztochen"
"Y20-64","BG4",2005,8.7,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2005,7.4,"Yugozapaden"
"Y20-64","BG42",2005,10.7,"Yuzhen tsentralen"
"Y20-64","CH",2005,4.3,"Switzerland"
"Y20-64","CH0",2005,4.3,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2005,6.2,"Région lémanique"
"Y20-64","CH02",2005,3.7,"Espace Mittelland"
"Y20-64","CH03",2005,3.9,"Nordwestschweiz"
"Y20-64","CH04",2005,4.2,"Zürich"
"Y20-64","CH05",2005,3.8,"Ostschweiz"
"Y20-64","CH06",2005,2.7,"Zentralschweiz"
"Y20-64","CH07",2005,5.8,"Ticino"
"Y20-64","CY",2005,5.2,"Cyprus"
"Y20-64","CY0",2005,5.2,"Kypros"
"Y20-64","CY00",2005,5.2,"Kypros"
"Y20-64","CZ",2005,7.6,"Czech Republic"
"Y20-64","CZ0",2005,7.6,"Ceská republika"
"Y20-64","CZ01",2005,3.5,"Praha"
"Y20-64","CZ02",2005,5,"Strední Cechy"
"Y20-64","CZ03",2005,4.8,"Jihozápad"
"Y20-64","CZ04",2005,12.5,"Severozápad"
"Y20-64","CZ05",2005,5.3,"Severovýchod"
"Y20-64","CZ06",2005,7.4,"Jihovýchod"
"Y20-64","CZ07",2005,9.4,"Strední Morava"
"Y20-64","CZ08",2005,13.3,"Moravskoslezsko"
"Y20-64","DE",2005,11.2,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2005,7,"Baden-Württemberg"
"Y20-64","DE11",2005,7.3,"Stuttgart"
"Y20-64","DE12",2005,7.5,"Karlsruhe"
"Y20-64","DE13",2005,6.2,"Freiburg"
"Y20-64","DE14",2005,6.8,"Tübingen"
"Y20-64","DE2",2005,6.9,"Bayern"
"Y20-64","DE21",2005,5.7,"Oberbayern"
"Y20-64","DE22",2005,6.3,"Niederbayern"
"Y20-64","DE23",2005,6.5,"Oberpfalz"
"Y20-64","DE24",2005,10,"Oberfranken"
"Y20-64","DE25",2005,8.6,"Mittelfranken"
"Y20-64","DE26",2005,7.9,"Unterfranken"
"Y20-64","DE27",2005,6.6,"Schwaben"
"Y20-64","DE3",2005,19.3,"Berlin"
"Y20-64","DE30",2005,19.3,"Berlin"
"Y20-64","DE4",2005,18.4,"Brandenburg"
"Y20-64","DE40",2005,18.4,"Brandenburg"
"Y20-64","DE5",2005,16.8,"Bremen"
"Y20-64","DE50",2005,16.8,"Bremen"
"Y20-64","DE6",2005,10.5,"Hamburg"
"Y20-64","DE60",2005,10.5,"Hamburg"
"Y20-64","DE7",2005,8.4,"Hessen"
"Y20-64","DE71",2005,8,"Darmstadt"
"Y20-64","DE72",2005,8.8,"Gießen"
"Y20-64","DE73",2005,9.3,"Kassel"
"Y20-64","DE8",2005,21.9,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2005,21.9,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2005,10.4,"Niedersachsen"
"Y20-64","DE91",2005,11.7,"Braunschweig"
"Y20-64","DE92",2005,10.2,"Hannover"
"Y20-64","DE93",2005,9.8,"Lüneburg"
"Y20-64","DE94",2005,10.2,"Weser-Ems"
"Y20-64","DEA",2005,10.4,"Nordrhein-Westfalen"
"Y20-64","DEA1",2005,10.6,"Düsseldorf"
"Y20-64","DEA2",2005,9.2,"Köln"
"Y20-64","DEA3",2005,9.5,"Münster"
"Y20-64","DEA4",2005,10.1,"Detmold"
"Y20-64","DEA5",2005,12.1,"Arnsberg"
"Y20-64","DEB",2005,8.7,"Rheinland-Pfalz"
"Y20-64","DEB1",2005,8.7,"Koblenz"
"Y20-64","DEB2",2005,7.4,"Trier"
"Y20-64","DEB3",2005,9.1,"Rheinhessen-Pfalz"
"Y20-64","DEC",2005,10.6,"Saarland"
"Y20-64","DEC0",2005,10.6,"Saarland"
"Y20-64","DED",2005,19,"Sachsen"
"Y20-64","DED2",2005,18.6,"Dresden"
"Y20-64","DED4",2005,18.5,"Chemnitz"
"Y20-64","DED5",2005,20.3,"Leipzig"
"Y20-64","DEE",2005,20.6,"Sachsen-Anhalt"
"Y20-64","DEE0",2005,20.6,"Sachsen-Anhalt"
"Y20-64","DEF",2005,10.2,"Schleswig-Holstein"
"Y20-64","DEF0",2005,10.2,"Schleswig-Holstein"
"Y20-64","DEG",2005,17.4,"Thüringen"
"Y20-64","DEG0",2005,17.4,"Thüringen"
"Y20-64","DK",2005,4.6,"Denmark"
"Y20-64","DK0",2005,4.6,"Danmark"
"Y20-64","EA17",2005,8.8,"Euro area (17 countries)"
"Y20-64","EA18",2005,8.8,"Euro area (18 countries)"
"Y20-64","EA19",2005,8.8,"Euro area (19 countries)"
"Y20-64","EE",2005,7.9,"Estonia"
"Y20-64","EE0",2005,7.9,"Eesti"
"Y20-64","EE00",2005,7.9,"Eesti"
"Y20-64","EL",2005,9.8,"Greece"
"Y20-64","EL1",2005,11.4,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2005,11.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2005,11,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2005,17.9,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2005,9.7,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2005,10,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2005,11.4,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2005,8.6,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2005,10.7,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2005,10.6,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2005,8.3,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2005,8.9,"Attiki"
"Y20-64","EL30",2005,8.9,"Attiki"
"Y20-64","EL4",2005,8.2,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2005,9.5,"Voreio Aigaio"
"Y20-64","EL42",2005,9.6,"Notio Aigaio"
"Y20-64","EL43",2005,7.1,"Kriti"
"Y20-64","ES",2005,8.7,"Spain"
"Y20-64","ES1",2005,9.5,"Noroeste (ES)"
"Y20-64","ES11",2005,9.7,"Galicia"
"Y20-64","ES12",2005,9.9,"Principado de Asturias"
"Y20-64","ES13",2005,8.2,"Cantabria"
"Y20-64","ES2",2005,6.4,"Noreste (ES)"
"Y20-64","ES21",2005,7.1,"País Vasco"
"Y20-64","ES22",2005,5.4,"Comunidad Foral de Navarra"
"Y20-64","ES23",2005,5.8,"La Rioja"
"Y20-64","ES24",2005,5.7,"Aragón"
"Y20-64","ES3",2005,6.4,"Comunidad de Madrid"
"Y20-64","ES30",2005,6.4,"Comunidad de Madrid"
"Y20-64","ES4",2005,9.8,"Centro (ES)"
"Y20-64","ES41",2005,8.5,"Castilla y León"
"Y20-64","ES42",2005,8.7,"Castilla-la Mancha"
"Y20-64","ES43",2005,14.9,"Extremadura"
"Y20-64","ES5",2005,7.1,"Este (ES)"
"Y20-64","ES51",2005,6.5,"Cataluña"
"Y20-64","ES52",2005,8.3,"Comunidad Valenciana"
"Y20-64","ES53",2005,6.2,"Illes Balears"
"Y20-64","ES6",2005,12.3,"Sur (ES)"
"Y20-64","ES61",2005,13.1,"Andalucía"
"Y20-64","ES62",2005,7.5,"Región de Murcia"
"Y20-64","ES63",2005,18.2,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2005,13.9,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2005,11,"Canarias (ES)"
"Y20-64","ES70",2005,11,"Canarias (ES)"
"Y20-64","EU15",2005,7.8,"European Union (15 countries)"
"Y20-64","EU27",2005,8.6,"European Union (27 countries)"
"Y20-64","EU28",2005,8.7,"European Union (28 countries)"
"Y20-64","FI",2005,7.7,"Finland"
"Y20-64","FI1",2005,7.7,"Manner-Suomi"
"Y20-64","FI19",2005,8.1,"Länsi-Suomi"
"Y20-64","FI1B",2005,5.4,"Helsinki-Uusimaa"
"Y20-64","FI1C",2005,7.4,"Etelä-Suomi"
"Y20-64","FI1D",2005,10.5,"Pohjois- ja Itä-Suomi"
"Y20-64","FI2",2005,NA,"Åland"
"Y20-64","FI20",2005,NA,"Åland"
"Y20-64","FR",2005,8.6,"France"
"Y20-64","FR1",2005,8.4,"Île de France"
"Y20-64","FR10",2005,8.4,"Île de France"
"Y20-64","FR2",2005,7.7,"Bassin Parisien"
"Y20-64","FR21",2005,9.3,"Champagne-Ardenne"
"Y20-64","FR22",2005,9.5,"Picardie"
"Y20-64","FR23",2005,7.3,"Haute-Normandie"
"Y20-64","FR24",2005,6.3,"Centre (FR)"
"Y20-64","FR25",2005,7.4,"Basse-Normandie"
"Y20-64","FR26",2005,6.9,"Bourgogne"
"Y20-64","FR3",2005,12,"Nord - Pas-de-Calais"
"Y20-64","FR30",2005,12,"Nord - Pas-de-Calais"
"Y20-64","FR4",2005,7.5,"Est (FR)"
"Y20-64","FR41",2005,9.4,"Lorraine"
"Y20-64","FR42",2005,6,"Alsace"
"Y20-64","FR43",2005,6.4,"Franche-Comté"
"Y20-64","FR5",2005,6.9,"Ouest (FR)"
"Y20-64","FR51",2005,6.7,"Pays de la Loire"
"Y20-64","FR52",2005,6.6,"Bretagne"
"Y20-64","FR53",2005,8,"Poitou-Charentes"
"Y20-64","FR6",2005,6.7,"Sud-Ouest (FR)"
"Y20-64","FR61",2005,7.1,"Aquitaine"
"Y20-64","FR62",2005,6.5,"Midi-Pyrénées"
"Y20-64","FR63",2005,6,"Limousin"
"Y20-64","FR7",2005,7.5,"Centre-Est (FR)"
"Y20-64","FR71",2005,7.6,"Rhône-Alpes"
"Y20-64","FR72",2005,6.9,"Auvergne"
"Y20-64","FR8",2005,10.2,"Méditerranée"
"Y20-64","FR81",2005,11.2,"Languedoc-Roussillon"
"Y20-64","FR82",2005,9.8,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2005,9.8,"Corse"
"Y20-64","FR9",2005,25.3,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2005,25.6,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2005,18.4,"Martinique (NUTS 2010)"
"Y20-64","FR93",2005,24.3,"Guyane (NUTS 2010)"
"Y20-64","FR94",2005,28.9,"Réunion (NUTS 2010)"
"Y20-64","HR",2005,12.2,"Croatia"
"Y20-64","HR0",2005,12.2,"Hrvatska"
"Y20-64","HU",2005,7,"Hungary"
"Y20-64","HU1",2005,5,"Közép-Magyarország"
"Y20-64","HU10",2005,5,"Közép-Magyarország"
"Y20-64","HU2",2005,6.6,"Dunántúl"
"Y20-64","HU21",2005,6.1,"Közép-Dunántúl"
"Y20-64","HU22",2005,5.8,"Nyugat-Dunántúl"
"Y20-64","HU23",2005,8.3,"Dél-Dunántúl"
"Y20-64","HU3",2005,8.9,"Alföld és Észak"
"Y20-64","HU31",2005,10.2,"Észak-Magyarország"
"Y20-64","HU32",2005,8.7,"Észak-Alföld"
"Y20-64","HU33",2005,7.9,"Dél-Alföld"
"Y20-64","IE",2005,4.1,"Ireland"
"Y20-64","IE0",2005,4.1,"Éire/Ireland"
"Y20-64","IE01",2005,4.2,"Border, Midland and Western"
"Y20-64","IE02",2005,4,"Southern and Eastern"
"Y20-64","IS",2005,2.1,"Iceland"
"Y20-64","IS0",2005,2.1,"Ísland"
"Y20-64","IS00",2005,2.1,"Ísland"
"Y20-64","IT",2005,7.4,"Italy"
"Y20-64","ITC",2005,4.1,"Nord-Ovest"
"Y20-64","ITC1",2005,4.4,"Piemonte"
"Y20-64","ITC2",2005,3.2,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2005,5.4,"Liguria"
"Y20-64","ITC4",2005,3.8,"Lombardia"
"Y20-64","ITF",2005,13.2,"Sud"
"Y20-64","ITF1",2005,7.6,"Abruzzo"
"Y20-64","ITF2",2005,9.3,"Molise"
"Y20-64","ITF3",2005,14.3,"Campania"
"Y20-64","ITF4",2005,13.9,"Puglia"
"Y20-64","ITF5",2005,11.9,"Basilicata"
"Y20-64","ITF6",2005,13.7,"Calabria"
"Y20-64","ITG",2005,14.5,"Isole"
"Y20-64","ITG1",2005,15.3,"Sicilia"
"Y20-64","ITG2",2005,12.5,"Sardegna"
"Y20-64","ITH",2005,3.8,"Nord-Est"
"Y20-64","ITH1",2005,2.5,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2005,3.4,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2005,4,"Veneto"
"Y20-64","ITH4",2005,4.1,"Friuli-Venezia Giulia"
"Y20-64","ITH5",2005,3.7,"Emilia-Romagna"
"Y20-64","ITI",2005,6.2,"Centro (IT)"
"Y20-64","ITI1",2005,5.2,"Toscana"
"Y20-64","ITI2",2005,5.6,"Umbria"
"Y20-64","ITI3",2005,4.7,"Marche"
"Y20-64","ITI4",2005,7.4,"Lazio"
"Y20-64","LT",2005,8.3,"Lithuania"
"Y20-64","LT0",2005,8.3,"Lietuva"
"Y20-64","LT00",2005,8.3,"Lietuva"
"Y20-64","LU",2005,4.3,"Luxembourg"
"Y20-64","LU0",2005,4.3,"Luxembourg"
"Y20-64","LU00",2005,4.3,"Luxembourg"
"Y20-64","LV",2005,9.7,"Latvia"
"Y20-64","LV0",2005,9.7,"Latvija"
"Y20-64","LV00",2005,9.7,"Latvija"
"Y20-64","MT",2005,5.6,"Malta"
"Y20-64","MT0",2005,5.6,"Malta"
"Y20-64","MT00",2005,5.6,"Malta"
"Y20-64","NL",2005,4.3,"Netherlands"
"Y20-64","NL1",2005,5.3,"Noord-Nederland"
"Y20-64","NL11",2005,6.3,"Groningen"
"Y20-64","NL12",2005,4.6,"Friesland (NL)"
"Y20-64","NL13",2005,5.2,"Drenthe"
"Y20-64","NL2",2005,4.3,"Oost-Nederland"
"Y20-64","NL21",2005,4.6,"Overijssel"
"Y20-64","NL22",2005,3.9,"Gelderland"
"Y20-64","NL23",2005,5.8,"Flevoland"
"Y20-64","NL3",2005,4.2,"West-Nederland"
"Y20-64","NL31",2005,3.3,"Utrecht"
"Y20-64","NL32",2005,4.6,"Noord-Holland"
"Y20-64","NL33",2005,4.4,"Zuid-Holland"
"Y20-64","NL34",2005,3.2,"Zeeland"
"Y20-64","NL4",2005,4.1,"Zuid-Nederland"
"Y20-64","NL41",2005,3.6,"Noord-Brabant"
"Y20-64","NL42",2005,5.1,"Limburg (NL)"
"Y20-64","NO",2005,3.8,"Norway"
"Y20-64","NO0",2005,3.8,"Norge"
"Y20-64","NO01",2005,4.2,"Oslo og Akershus"
"Y20-64","NO02",2005,3.5,"Hedmark og Oppland"
"Y20-64","NO03",2005,4.1,"Sør-Østlandet"
"Y20-64","NO04",2005,3.6,"Agder og Rogaland"
"Y20-64","NO05",2005,3.4,"Vestlandet"
"Y20-64","NO06",2005,2.9,"Trøndelag"
"Y20-64","NO07",2005,4.2,"Nord-Norge"
"Y20-64","PL",2005,17.7,"Poland"
"Y20-64","PL1",2005,15.9,"Region Centralny"
"Y20-64","PL11",2005,17.4,"Lódzkie"
"Y20-64","PL12",2005,14.9,"Mazowieckie"
"Y20-64","PL2",2005,17.4,"Region Poludniowy"
"Y20-64","PL21",2005,15.5,"Malopolskie"
"Y20-64","PL22",2005,18.6,"Slaskie"
"Y20-64","PL3",2005,16.3,"Region Wschodni"
"Y20-64","PL31",2005,14.6,"Lubelskie"
"Y20-64","PL32",2005,17,"Podkarpackie"
"Y20-64","PL33",2005,19.4,"Swietokrzyskie"
"Y20-64","PL34",2005,14.5,"Podlaskie"
"Y20-64","PL4",2005,18.7,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2005,16.9,"Wielkopolskie"
"Y20-64","PL42",2005,22.3,"Zachodniopomorskie"
"Y20-64","PL43",2005,18.9,"Lubuskie"
"Y20-64","PL5",2005,21.2,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2005,22.5,"Dolnoslaskie"
"Y20-64","PL52",2005,17,"Opolskie"
"Y20-64","PL6",2005,19.4,"Region Pólnocny"
"Y20-64","PL61",2005,19.7,"Kujawsko-Pomorskie"
"Y20-64","PL62",2005,20.2,"Warminsko-Mazurskie"
"Y20-64","PL63",2005,18.6,"Pomorskie"
"Y20-64","PT",2005,7.8,"Portugal"
"Y20-64","PT1",2005,7.9,"Continente"
"Y20-64","PT11",2005,9,"Norte"
"Y20-64","PT15",2005,6.1,"Algarve"
"Y20-64","PT16",2005,5.7,"Centro (PT)"
"Y20-64","PT17",2005,8.5,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2005,9,"Alentejo"
"Y20-64","PT2",2005,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2005,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2005,4.4,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2005,4.4,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2005,7,"Romania"
"Y20-64","RO1",2005,6.8,"Macroregiunea unu"
"Y20-64","RO11",2005,5.6,"Nord-Vest"
"Y20-64","RO12",2005,8,"Centru"
"Y20-64","RO2",2005,6.5,"Macroregiunea doi"
"Y20-64","RO21",2005,5.7,"Nord-Est"
"Y20-64","RO22",2005,7.6,"Sud-Est"
"Y20-64","RO3",2005,8,"Macroregiunea trei"
"Y20-64","RO31",2005,9.2,"Sud - Muntenia"
"Y20-64","RO32",2005,6.4,"Bucuresti - Ilfov"
"Y20-64","RO4",2005,6.7,"Macroregiunea patru"
"Y20-64","RO41",2005,7,"Sud-Vest Oltenia"
"Y20-64","RO42",2005,6.5,"Vest"
"Y20-64","SE",2005,6.8,"Sweden"
"Y20-64","SE1",2005,6.5,"Östra Sverige"
"Y20-64","SE11",2005,5.9,"Stockholm"
"Y20-64","SE12",2005,7.3,"Östra Mellansverige"
"Y20-64","SE2",2005,6.7,"Södra Sverige"
"Y20-64","SE21",2005,5.4,"Småland med öarna"
"Y20-64","SE22",2005,8.1,"Sydsverige"
"Y20-64","SE23",2005,6.3,"Västsverige"
"Y20-64","SE3",2005,7.9,"Norra Sverige"
"Y20-64","SE31",2005,8.2,"Norra Mellansverige"
"Y20-64","SE32",2005,7.6,"Mellersta Norrland"
"Y20-64","SE33",2005,7.7,"Övre Norrland"
"Y20-64","SI",2005,6.5,"Slovenia"
"Y20-64","SI0",2005,6.5,"Slovenija"
"Y20-64","SI01",2005,7.5,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2005,5.2,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2005,15.7,"Slovakia"
"Y20-64","SK0",2005,15.7,"Slovensko"
"Y20-64","SK01",2005,5.1,"Bratislavský kraj"
"Y20-64","SK02",2005,12.2,"Západné Slovensko"
"Y20-64","SK03",2005,18.9,"Stredné Slovensko"
"Y20-64","SK04",2005,22,"Východné Slovensko"
"Y20-64","UK",2005,4,"United Kingdom"
"Y20-64","UKC",2005,4.9,"North East (UK)"
"Y20-64","UKC1",2005,4.6,"Tees Valley and Durham"
"Y20-64","UKC2",2005,5.2,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2005,3.7,"North West (UK)"
"Y20-64","UKD1",2005,3.1,"Cumbria"
"Y20-64","UKD3",2005,3.9,"Greater Manchester"
"Y20-64","UKD4",2005,3.4,"Lancashire"
"Y20-64","UKD6",2005,2.5,"Cheshire"
"Y20-64","UKD7",2005,4.5,"Merseyside"
"Y20-64","UKE",2005,3.8,"Yorkshire and The Humber"
"Y20-64","UKE1",2005,4.4,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2005,2.3,"North Yorkshire"
"Y20-64","UKE3",2005,4.5,"South Yorkshire"
"Y20-64","UKE4",2005,3.7,"West Yorkshire"
"Y20-64","UKF",2005,3.5,"East Midlands (UK)"
"Y20-64","UKF1",2005,3.5,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2005,3.6,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2005,3,"Lincolnshire"
"Y20-64","UKG",2005,3.9,"West Midlands (UK)"
"Y20-64","UKG1",2005,2.2,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2005,3.2,"Shropshire and Staffordshire"
"Y20-64","UKG3",2005,5.3,"West Midlands"
"Y20-64","UKH",2005,3.3,"East of England"
"Y20-64","UKH1",2005,3.4,"East Anglia"
"Y20-64","UKH2",2005,3.3,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2005,3.1,"Essex"
"Y20-64","UKI",2005,6.2,"London"
"Y20-64","UKI1",2005,7.1,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2005,5.6,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2005,3.2,"South East (UK)"
"Y20-64","UKJ1",2005,2.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2005,3.2,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2005,3.5,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2005,3.6,"Kent"
"Y20-64","UKK",2005,3,"South West (UK)"
"Y20-64","UKK1",2005,2.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2005,3.1,"Dorset and Somerset"
"Y20-64","UKK3",2005,2.8,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2005,3.1,"Devon"
"Y20-64","UKL",2005,3.4,"Wales"
"Y20-64","UKL1",2005,3.9,"West Wales and The Valleys"
"Y20-64","UKL2",2005,2.7,"East Wales"
"Y20-64","UKM",2005,4.4,"Scotland"
"Y20-64","UKM2",2005,4.5,"Eastern Scotland"
"Y20-64","UKM3",2005,4.9,"South Western Scotland"
"Y20-64","UKM5",2005,3.3,"North Eastern Scotland"
"Y20-64","UKM6",2005,3,"Highlands and Islands"
"Y20-64","UKN",2005,4.1,"Northern Ireland (UK)"
"Y20-64","UKN0",2005,4.1,"Northern Ireland (UK)"
"Y_GE15","AT",2005,5.6,"Austria"
"Y_GE15","AT1",2005,7.3,"Ostösterreich"
"Y_GE15","AT11",2005,5.8,"Burgenland (AT)"
"Y_GE15","AT12",2005,4.7,"Niederösterreich"
"Y_GE15","AT13",2005,9.9,"Wien"
"Y_GE15","AT2",2005,4.8,"Südösterreich"
"Y_GE15","AT21",2005,5.3,"Kärnten"
"Y_GE15","AT22",2005,4.5,"Steiermark"
"Y_GE15","AT3",2005,4.3,"Westösterreich"
"Y_GE15","AT31",2005,4.4,"Oberösterreich"
"Y_GE15","AT32",2005,3.6,"Salzburg"
"Y_GE15","AT33",2005,3.9,"Tirol"
"Y_GE15","AT34",2005,5.5,"Vorarlberg"
"Y_GE15","BE",2005,8.4,"Belgium"
"Y_GE15","BE1",2005,16.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2005,16.3,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2005,5.4,"Vlaams Gewest"
"Y_GE15","BE21",2005,6.2,"Prov. Antwerpen"
"Y_GE15","BE22",2005,7.1,"Prov. Limburg (BE)"
"Y_GE15","BE23",2005,4.9,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2005,4.4,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2005,4.7,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2005,11.8,"Région wallonne"
"Y_GE15","BE31",2005,9,"Prov. Brabant Wallon"
"Y_GE15","BE32",2005,14,"Prov. Hainaut"
"Y_GE15","BE33",2005,11.9,"Prov. Liège"
"Y_GE15","BE34",2005,7.9,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2005,10.4,"Prov. Namur"
"Y_GE15","BG",2005,10.1,"Bulgaria"
"Y_GE15","BG3",2005,11.2,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2005,12.6,"Severozapaden"
"Y_GE15","BG32",2005,12.5,"Severen tsentralen"
"Y_GE15","BG33",2005,12.1,"Severoiztochen"
"Y_GE15","BG34",2005,8.3,"Yugoiztochen"
"Y_GE15","BG4",2005,8.9,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2005,7.6,"Yugozapaden"
"Y_GE15","BG42",2005,11,"Yuzhen tsentralen"
"Y_GE15","CH",2005,4.4,"Switzerland"
"Y_GE15","CH0",2005,4.4,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2005,6.5,"Région lémanique"
"Y_GE15","CH02",2005,4,"Espace Mittelland"
"Y_GE15","CH03",2005,4.1,"Nordwestschweiz"
"Y_GE15","CH04",2005,4.2,"Zürich"
"Y_GE15","CH05",2005,3.8,"Ostschweiz"
"Y_GE15","CH06",2005,2.9,"Zentralschweiz"
"Y_GE15","CH07",2005,6.1,"Ticino"
"Y_GE15","CY",2005,5.3,"Cyprus"
"Y_GE15","CY0",2005,5.3,"Kypros"
"Y_GE15","CY00",2005,5.3,"Kypros"
"Y_GE15","CZ",2005,7.9,"Czech Republic"
"Y_GE15","CZ0",2005,7.9,"Ceská republika"
"Y_GE15","CZ01",2005,3.5,"Praha"
"Y_GE15","CZ02",2005,5.2,"Strední Cechy"
"Y_GE15","CZ03",2005,5.1,"Jihozápad"
"Y_GE15","CZ04",2005,13.5,"Severozápad"
"Y_GE15","CZ05",2005,5.6,"Severovýchod"
"Y_GE15","CZ06",2005,7.7,"Jihovýchod"
"Y_GE15","CZ07",2005,9.7,"Strední Morava"
"Y_GE15","CZ08",2005,13.9,"Moravskoslezsko"
"Y_GE15","DE",2005,11.2,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2005,7.1,"Baden-Württemberg"
"Y_GE15","DE11",2005,7.3,"Stuttgart"
"Y_GE15","DE12",2005,7.6,"Karlsruhe"
"Y_GE15","DE13",2005,6.4,"Freiburg"
"Y_GE15","DE14",2005,6.8,"Tübingen"
"Y_GE15","DE2",2005,7.1,"Bayern"
"Y_GE15","DE21",2005,5.8,"Oberbayern"
"Y_GE15","DE22",2005,6.4,"Niederbayern"
"Y_GE15","DE23",2005,6.5,"Oberpfalz"
"Y_GE15","DE24",2005,10.3,"Oberfranken"
"Y_GE15","DE25",2005,8.7,"Mittelfranken"
"Y_GE15","DE26",2005,8.2,"Unterfranken"
"Y_GE15","DE27",2005,6.5,"Schwaben"
"Y_GE15","DE3",2005,19.3,"Berlin"
"Y_GE15","DE30",2005,19.3,"Berlin"
"Y_GE15","DE4",2005,18.2,"Brandenburg"
"Y_GE15","DE40",2005,18.2,"Brandenburg"
"Y_GE15","DE5",2005,16.7,"Bremen"
"Y_GE15","DE50",2005,16.7,"Bremen"
"Y_GE15","DE6",2005,10.5,"Hamburg"
"Y_GE15","DE60",2005,10.5,"Hamburg"
"Y_GE15","DE7",2005,8.5,"Hessen"
"Y_GE15","DE71",2005,8.1,"Darmstadt"
"Y_GE15","DE72",2005,9,"Gießen"
"Y_GE15","DE73",2005,9.3,"Kassel"
"Y_GE15","DE8",2005,21.4,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2005,21.4,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2005,10.4,"Niedersachsen"
"Y_GE15","DE91",2005,11.6,"Braunschweig"
"Y_GE15","DE92",2005,10.5,"Hannover"
"Y_GE15","DE93",2005,9.7,"Lüneburg"
"Y_GE15","DE94",2005,10.2,"Weser-Ems"
"Y_GE15","DEA",2005,10.5,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2005,10.6,"Düsseldorf"
"Y_GE15","DEA2",2005,9.4,"Köln"
"Y_GE15","DEA3",2005,9.5,"Münster"
"Y_GE15","DEA4",2005,10.2,"Detmold"
"Y_GE15","DEA5",2005,12.2,"Arnsberg"
"Y_GE15","DEB",2005,8.8,"Rheinland-Pfalz"
"Y_GE15","DEB1",2005,8.7,"Koblenz"
"Y_GE15","DEB2",2005,7.3,"Trier"
"Y_GE15","DEB3",2005,9.2,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2005,10.8,"Saarland"
"Y_GE15","DEC0",2005,10.8,"Saarland"
"Y_GE15","DED",2005,18.7,"Sachsen"
"Y_GE15","DED2",2005,18.3,"Dresden"
"Y_GE15","DED4",2005,18,"Chemnitz"
"Y_GE15","DED5",2005,20.3,"Leipzig"
"Y_GE15","DEE",2005,20.4,"Sachsen-Anhalt"
"Y_GE15","DEE0",2005,20.4,"Sachsen-Anhalt"
"Y_GE15","DEF",2005,10.3,"Schleswig-Holstein"
"Y_GE15","DEF0",2005,10.3,"Schleswig-Holstein"
"Y_GE15","DEG",2005,17.2,"Thüringen"
"Y_GE15","DEG0",2005,17.2,"Thüringen"
"Y_GE15","DK",2005,4.8,"Denmark"
"Y_GE15","DK0",2005,4.8,"Danmark"
"Y_GE15","EA17",2005,9,"Euro area (17 countries)"
"Y_GE15","EA18",2005,9,"Euro area (18 countries)"
"Y_GE15","EA19",2005,9,"Euro area (19 countries)"
"Y_GE15","EE",2005,8,"Estonia"
"Y_GE15","EE0",2005,8,"Eesti"
"Y_GE15","EE00",2005,8,"Eesti"
"Y_GE15","EL",2005,10,"Greece"
"Y_GE15","EL1",2005,11.5,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2005,11.9,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2005,11.2,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2005,18.1,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2005,9.4,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2005,10.2,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2005,11.5,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2005,8.6,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2005,10.7,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2005,11,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2005,8.6,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2005,9.1,"Attiki"
"Y_GE15","EL30",2005,9.1,"Attiki"
"Y_GE15","EL4",2005,8.4,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2005,10.6,"Voreio Aigaio"
"Y_GE15","EL42",2005,9.5,"Notio Aigaio"
"Y_GE15","EL43",2005,7.2,"Kriti"
"Y_GE15","ES",2005,9.1,"Spain"
"Y_GE15","ES1",2005,9.7,"Noroeste (ES)"
"Y_GE15","ES11",2005,9.9,"Galicia"
"Y_GE15","ES12",2005,10,"Principado de Asturias"
"Y_GE15","ES13",2005,8.5,"Cantabria"
"Y_GE15","ES2",2005,6.6,"Noreste (ES)"
"Y_GE15","ES21",2005,7.4,"País Vasco"
"Y_GE15","ES22",2005,5.7,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2005,6.4,"La Rioja"
"Y_GE15","ES24",2005,5.9,"Aragón"
"Y_GE15","ES3",2005,6.8,"Comunidad de Madrid"
"Y_GE15","ES30",2005,6.8,"Comunidad de Madrid"
"Y_GE15","ES4",2005,10.2,"Centro (ES)"
"Y_GE15","ES41",2005,8.7,"Castilla y León"
"Y_GE15","ES42",2005,9.2,"Castilla-la Mancha"
"Y_GE15","ES43",2005,15.7,"Extremadura"
"Y_GE15","ES5",2005,7.6,"Este (ES)"
"Y_GE15","ES51",2005,6.9,"Cataluña"
"Y_GE15","ES52",2005,8.9,"Comunidad Valenciana"
"Y_GE15","ES53",2005,7.2,"Illes Balears"
"Y_GE15","ES6",2005,13,"Sur (ES)"
"Y_GE15","ES61",2005,13.8,"Andalucía"
"Y_GE15","ES62",2005,8,"Región de Murcia"
"Y_GE15","ES63",2005,19.4,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2005,14.3,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2005,11.7,"Canarias (ES)"
"Y_GE15","ES70",2005,11.7,"Canarias (ES)"
"Y_GE15","EU15",2005,8.2,"European Union (15 countries)"
"Y_GE15","EU27",2005,8.9,"European Union (27 countries)"
"Y_GE15","EU28",2005,9,"European Union (28 countries)"
"Y_GE15","FI",2005,8.4,"Finland"
"Y_GE15","FI1",2005,8.4,"Manner-Suomi"
"Y_GE15","FI19",2005,8.8,"Länsi-Suomi"
"Y_GE15","FI1B",2005,6.1,"Helsinki-Uusimaa"
"Y_GE15","FI1C",2005,8.1,"Etelä-Suomi"
"Y_GE15","FI1D",2005,11.4,"Pohjois- ja Itä-Suomi"
"Y_GE15","FI2",2005,NA,"Åland"
"Y_GE15","FI20",2005,NA,"Åland"
"Y_GE15","FR",2005,8.9,"France"
"Y_GE15","FR1",2005,8.6,"Île de France"
"Y_GE15","FR10",2005,8.6,"Île de France"
"Y_GE15","FR2",2005,8.1,"Bassin Parisien"
"Y_GE15","FR21",2005,9.7,"Champagne-Ardenne"
"Y_GE15","FR22",2005,10.2,"Picardie"
"Y_GE15","FR23",2005,7.7,"Haute-Normandie"
"Y_GE15","FR24",2005,6.9,"Centre (FR)"
"Y_GE15","FR25",2005,7.7,"Basse-Normandie"
"Y_GE15","FR26",2005,7.2,"Bourgogne"
"Y_GE15","FR3",2005,12.8,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2005,12.8,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2005,8.2,"Est (FR)"
"Y_GE15","FR41",2005,9.9,"Lorraine"
"Y_GE15","FR42",2005,6.9,"Alsace"
"Y_GE15","FR43",2005,7,"Franche-Comté"
"Y_GE15","FR5",2005,7.3,"Ouest (FR)"
"Y_GE15","FR51",2005,7.2,"Pays de la Loire"
"Y_GE15","FR52",2005,6.7,"Bretagne"
"Y_GE15","FR53",2005,8.4,"Poitou-Charentes"
"Y_GE15","FR6",2005,6.9,"Sud-Ouest (FR)"
"Y_GE15","FR61",2005,7.3,"Aquitaine"
"Y_GE15","FR62",2005,6.7,"Midi-Pyrénées"
"Y_GE15","FR63",2005,6.3,"Limousin"
"Y_GE15","FR7",2005,7.7,"Centre-Est (FR)"
"Y_GE15","FR71",2005,7.8,"Rhône-Alpes"
"Y_GE15","FR72",2005,7.1,"Auvergne"
"Y_GE15","FR8",2005,10.5,"Méditerranée"
"Y_GE15","FR81",2005,11.5,"Languedoc-Roussillon"
"Y_GE15","FR82",2005,10.1,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2005,10.2,"Corse"
"Y_GE15","FR9",2005,26.1,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2005,25.9,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2005,18.7,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2005,24.8,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2005,30.1,"Réunion (NUTS 2010)"
"Y_GE15","HR",2005,12.6,"Croatia"
"Y_GE15","HR0",2005,12.6,"Hrvatska"
"Y_GE15","HU",2005,7.2,"Hungary"
"Y_GE15","HU1",2005,5.1,"Közép-Magyarország"
"Y_GE15","HU10",2005,5.1,"Közép-Magyarország"
"Y_GE15","HU2",2005,6.9,"Dunántúl"
"Y_GE15","HU21",2005,6.3,"Közép-Dunántúl"
"Y_GE15","HU22",2005,5.9,"Nyugat-Dunántúl"
"Y_GE15","HU23",2005,8.8,"Dél-Dunántúl"
"Y_GE15","HU3",2005,9.2,"Alföld és Észak"
"Y_GE15","HU31",2005,10.6,"Észak-Magyarország"
"Y_GE15","HU32",2005,9,"Észak-Alföld"
"Y_GE15","HU33",2005,8.1,"Dél-Alföld"
"Y_GE15","IE",2005,4.3,"Ireland"
"Y_GE15","IE0",2005,4.3,"Éire/Ireland"
"Y_GE15","IE01",2005,4.4,"Border, Midland and Western"
"Y_GE15","IE02",2005,4.3,"Southern and Eastern"
"Y_GE15","IS",2005,2.5,"Iceland"
"Y_GE15","IS0",2005,2.5,"Ísland"
"Y_GE15","IS00",2005,2.5,"Ísland"
"Y_GE15","IT",2005,7.7,"Italy"
"Y_GE15","ITC",2005,4.4,"Nord-Ovest"
"Y_GE15","ITC1",2005,4.7,"Piemonte"
"Y_GE15","ITC2",2005,3.2,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2005,5.8,"Liguria"
"Y_GE15","ITC4",2005,4.1,"Lombardia"
"Y_GE15","ITF",2005,13.7,"Sud"
"Y_GE15","ITF1",2005,7.9,"Abruzzo"
"Y_GE15","ITF2",2005,9.9,"Molise"
"Y_GE15","ITF3",2005,14.9,"Campania"
"Y_GE15","ITF4",2005,14.6,"Puglia"
"Y_GE15","ITF5",2005,12.3,"Basilicata"
"Y_GE15","ITF6",2005,14.2,"Calabria"
"Y_GE15","ITG",2005,15.2,"Isole"
"Y_GE15","ITG1",2005,16.1,"Sicilia"
"Y_GE15","ITG2",2005,12.8,"Sardegna"
"Y_GE15","ITH",2005,4,"Nord-Est"
"Y_GE15","ITH1",2005,2.7,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2005,3.6,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2005,4.2,"Veneto"
"Y_GE15","ITH4",2005,4.2,"Friuli-Venezia Giulia"
"Y_GE15","ITH5",2005,3.9,"Emilia-Romagna"
"Y_GE15","ITI",2005,6.4,"Centro (IT)"
"Y_GE15","ITI1",2005,5.4,"Toscana"
"Y_GE15","ITI2",2005,6,"Umbria"
"Y_GE15","ITI3",2005,4.9,"Marche"
"Y_GE15","ITI4",2005,7.7,"Lazio"
"Y_GE15","LT",2005,8.3,"Lithuania"
"Y_GE15","LT0",2005,8.3,"Lietuva"
"Y_GE15","LT00",2005,8.3,"Lietuva"
"Y_GE15","LU",2005,4.5,"Luxembourg"
"Y_GE15","LU0",2005,4.5,"Luxembourg"
"Y_GE15","LU00",2005,4.5,"Luxembourg"
"Y_GE15","LV",2005,10,"Latvia"
"Y_GE15","LV0",2005,10,"Latvija"
"Y_GE15","LV00",2005,10,"Latvija"
"Y_GE15","MT",2005,6.9,"Malta"
"Y_GE15","MT0",2005,6.9,"Malta"
"Y_GE15","MT00",2005,6.9,"Malta"
"Y_GE15","NL",2005,4.7,"Netherlands"
"Y_GE15","NL1",2005,5.7,"Noord-Nederland"
"Y_GE15","NL11",2005,6.6,"Groningen"
"Y_GE15","NL12",2005,4.9,"Friesland (NL)"
"Y_GE15","NL13",2005,5.7,"Drenthe"
"Y_GE15","NL2",2005,4.8,"Oost-Nederland"
"Y_GE15","NL21",2005,4.9,"Overijssel"
"Y_GE15","NL22",2005,4.3,"Gelderland"
"Y_GE15","NL23",2005,6.6,"Flevoland"
"Y_GE15","NL3",2005,4.7,"West-Nederland"
"Y_GE15","NL31",2005,3.8,"Utrecht"
"Y_GE15","NL32",2005,4.9,"Noord-Holland"
"Y_GE15","NL33",2005,4.9,"Zuid-Holland"
"Y_GE15","NL34",2005,3.3,"Zeeland"
"Y_GE15","NL4",2005,4.4,"Zuid-Nederland"
"Y_GE15","NL41",2005,3.9,"Noord-Brabant"
"Y_GE15","NL42",2005,5.4,"Limburg (NL)"
"Y_GE15","NO",2005,4.4,"Norway"
"Y_GE15","NO0",2005,4.4,"Norge"
"Y_GE15","NO01",2005,4.6,"Oslo og Akershus"
"Y_GE15","NO02",2005,4.2,"Hedmark og Oppland"
"Y_GE15","NO03",2005,4.7,"Sør-Østlandet"
"Y_GE15","NO04",2005,4.1,"Agder og Rogaland"
"Y_GE15","NO05",2005,4.1,"Vestlandet"
"Y_GE15","NO06",2005,3.5,"Trøndelag"
"Y_GE15","NO07",2005,5.1,"Nord-Norge"
"Y_GE15","PL",2005,17.7,"Poland"
"Y_GE15","PL1",2005,15.7,"Region Centralny"
"Y_GE15","PL11",2005,17.4,"Lódzkie"
"Y_GE15","PL12",2005,14.8,"Mazowieckie"
"Y_GE15","PL2",2005,17.4,"Region Poludniowy"
"Y_GE15","PL21",2005,15.3,"Malopolskie"
"Y_GE15","PL22",2005,19,"Slaskie"
"Y_GE15","PL3",2005,15.9,"Region Wschodni"
"Y_GE15","PL31",2005,14.3,"Lubelskie"
"Y_GE15","PL32",2005,16.7,"Podkarpackie"
"Y_GE15","PL33",2005,19,"Swietokrzyskie"
"Y_GE15","PL34",2005,14.4,"Podlaskie"
"Y_GE15","PL4",2005,18.9,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2005,17.2,"Wielkopolskie"
"Y_GE15","PL42",2005,22.7,"Zachodniopomorskie"
"Y_GE15","PL43",2005,19.1,"Lubuskie"
"Y_GE15","PL5",2005,21.4,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2005,22.8,"Dolnoslaskie"
"Y_GE15","PL52",2005,16.9,"Opolskie"
"Y_GE15","PL6",2005,19.7,"Region Pólnocny"
"Y_GE15","PL61",2005,19.8,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2005,20.4,"Warminsko-Mazurskie"
"Y_GE15","PL63",2005,18.9,"Pomorskie"
"Y_GE15","PT",2005,7.6,"Portugal"
"Y_GE15","PT1",2005,7.7,"Continente"
"Y_GE15","PT11",2005,8.8,"Norte"
"Y_GE15","PT15",2005,6.2,"Algarve"
"Y_GE15","PT16",2005,5.1,"Centro (PT)"
"Y_GE15","PT17",2005,8.6,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2005,9.1,"Alentejo"
"Y_GE15","PT2",2005,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2005,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2005,4.5,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2005,4.5,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2005,7.2,"Romania"
"Y_GE15","RO1",2005,7.1,"Macroregiunea unu"
"Y_GE15","RO11",2005,5.9,"Nord-Vest"
"Y_GE15","RO12",2005,8.4,"Centru"
"Y_GE15","RO2",2005,6.6,"Macroregiunea doi"
"Y_GE15","RO21",2005,5.7,"Nord-Est"
"Y_GE15","RO22",2005,7.9,"Sud-Est"
"Y_GE15","RO3",2005,8.3,"Macroregiunea trei"
"Y_GE15","RO31",2005,9.2,"Sud - Muntenia"
"Y_GE15","RO32",2005,6.9,"Bucuresti - Ilfov"
"Y_GE15","RO4",2005,6.6,"Macroregiunea patru"
"Y_GE15","RO41",2005,6.6,"Sud-Vest Oltenia"
"Y_GE15","RO42",2005,6.7,"Vest"
"Y_GE15","SE",2005,7.8,"Sweden"
"Y_GE15","SE1",2005,7.5,"Östra Sverige"
"Y_GE15","SE11",2005,6.9,"Stockholm"
"Y_GE15","SE12",2005,8.1,"Östra Mellansverige"
"Y_GE15","SE2",2005,7.6,"Södra Sverige"
"Y_GE15","SE21",2005,6.1,"Småland med öarna"
"Y_GE15","SE22",2005,8.9,"Sydsverige"
"Y_GE15","SE23",2005,7.4,"Västsverige"
"Y_GE15","SE3",2005,9,"Norra Sverige"
"Y_GE15","SE31",2005,9.2,"Norra Mellansverige"
"Y_GE15","SE32",2005,8.9,"Mellersta Norrland"
"Y_GE15","SE33",2005,8.8,"Övre Norrland"
"Y_GE15","SI",2005,6.5,"Slovenia"
"Y_GE15","SI0",2005,6.5,"Slovenija"
"Y_GE15","SI01",2005,7.6,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2005,5.2,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2005,16.3,"Slovakia"
"Y_GE15","SK0",2005,16.3,"Slovensko"
"Y_GE15","SK01",2005,5.3,"Bratislavský kraj"
"Y_GE15","SK02",2005,12.5,"Západné Slovensko"
"Y_GE15","SK03",2005,19.6,"Stredné Slovensko"
"Y_GE15","SK04",2005,23.1,"Východné Slovensko"
"Y_GE15","UK",2005,4.8,"United Kingdom"
"Y_GE15","UKC",2005,6.1,"North East (UK)"
"Y_GE15","UKC1",2005,5.9,"Tees Valley and Durham"
"Y_GE15","UKC2",2005,6.2,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2005,4.6,"North West (UK)"
"Y_GE15","UKD1",2005,3.8,"Cumbria"
"Y_GE15","UKD3",2005,4.9,"Greater Manchester"
"Y_GE15","UKD4",2005,4.3,"Lancashire"
"Y_GE15","UKD6",2005,3.2,"Cheshire"
"Y_GE15","UKD7",2005,5.6,"Merseyside"
"Y_GE15","UKE",2005,4.7,"Yorkshire and The Humber"
"Y_GE15","UKE1",2005,5.4,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2005,2.9,"North Yorkshire"
"Y_GE15","UKE3",2005,5.4,"South Yorkshire"
"Y_GE15","UKE4",2005,4.6,"West Yorkshire"
"Y_GE15","UKF",2005,4.3,"East Midlands (UK)"
"Y_GE15","UKF1",2005,4.3,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2005,4.6,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2005,3.7,"Lincolnshire"
"Y_GE15","UKG",2005,4.7,"West Midlands (UK)"
"Y_GE15","UKG1",2005,2.6,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2005,3.7,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2005,6.4,"West Midlands"
"Y_GE15","UKH",2005,3.9,"East of England"
"Y_GE15","UKH1",2005,4.1,"East Anglia"
"Y_GE15","UKH2",2005,3.8,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2005,3.8,"Essex"
"Y_GE15","UKI",2005,7,"London"
"Y_GE15","UKI1",2005,7.9,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2005,6.5,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2005,3.8,"South East (UK)"
"Y_GE15","UKJ1",2005,3.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2005,3.7,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2005,3.9,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2005,4.2,"Kent"
"Y_GE15","UKK",2005,3.6,"South West (UK)"
"Y_GE15","UKK1",2005,3.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2005,3.5,"Dorset and Somerset"
"Y_GE15","UKK3",2005,3.4,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2005,3.9,"Devon"
"Y_GE15","UKL",2005,4.5,"Wales"
"Y_GE15","UKL1",2005,5,"West Wales and The Valleys"
"Y_GE15","UKL2",2005,3.5,"East Wales"
"Y_GE15","UKM",2005,5.3,"Scotland"
"Y_GE15","UKM2",2005,5.1,"Eastern Scotland"
"Y_GE15","UKM3",2005,6.2,"South Western Scotland"
"Y_GE15","UKM5",2005,3.9,"North Eastern Scotland"
"Y_GE15","UKM6",2005,3.5,"Highlands and Islands"
"Y_GE15","UKN",2005,4.7,"Northern Ireland (UK)"
"Y_GE15","UKN0",2005,4.7,"Northern Ireland (UK)"
"Y_GE25","AT",2005,4.7,"Austria"
"Y_GE25","AT1",2005,6.1,"Ostösterreich"
"Y_GE25","AT11",2005,4.7,"Burgenland (AT)"
"Y_GE25","AT12",2005,4,"Niederösterreich"
"Y_GE25","AT13",2005,8.4,"Wien"
"Y_GE25","AT2",2005,3.9,"Südösterreich"
"Y_GE25","AT21",2005,4.3,"Kärnten"
"Y_GE25","AT22",2005,3.8,"Steiermark"
"Y_GE25","AT3",2005,3.5,"Westösterreich"
"Y_GE25","AT31",2005,3.8,"Oberösterreich"
"Y_GE25","AT32",2005,2.8,"Salzburg"
"Y_GE25","AT33",2005,3,"Tirol"
"Y_GE25","AT34",2005,4.5,"Vorarlberg"
"Y_GE25","BE",2005,7.1,"Belgium"
"Y_GE25","BE1",2005,14.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2005,14.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2005,4.5,"Vlaams Gewest"
"Y_GE25","BE21",2005,5.6,"Prov. Antwerpen"
"Y_GE25","BE22",2005,6,"Prov. Limburg (BE)"
"Y_GE25","BE23",2005,3.7,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2005,3.4,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2005,3.9,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2005,9.6,"Région wallonne"
"Y_GE25","BE31",2005,7.4,"Prov. Brabant Wallon"
"Y_GE25","BE32",2005,11.3,"Prov. Hainaut"
"Y_GE25","BE33",2005,10.3,"Prov. Liège"
"Y_GE25","BE34",2005,6,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2005,8,"Prov. Namur"
"Y_GE25","BG",2005,8.9,"Bulgaria"
"Y_GE25","BG3",2005,9.9,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2005,11,"Severozapaden"
"Y_GE25","BG32",2005,11.2,"Severen tsentralen"
"Y_GE25","BG33",2005,10.7,"Severoiztochen"
"Y_GE25","BG34",2005,7.2,"Yugoiztochen"
"Y_GE25","BG4",2005,7.9,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2005,6.9,"Yugozapaden"
"Y_GE25","BG42",2005,9.4,"Yuzhen tsentralen"
"Y_GE25","CH",2005,3.7,"Switzerland"
"Y_GE25","CH0",2005,3.7,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2005,5.5,"Région lémanique"
"Y_GE25","CH02",2005,3.3,"Espace Mittelland"
"Y_GE25","CH03",2005,3.6,"Nordwestschweiz"
"Y_GE25","CH04",2005,3.8,"Zürich"
"Y_GE25","CH05",2005,2.9,"Ostschweiz"
"Y_GE25","CH06",2005,2.4,"Zentralschweiz"
"Y_GE25","CH07",2005,4.9,"Ticino"
"Y_GE25","CY",2005,4.3,"Cyprus"
"Y_GE25","CY0",2005,4.3,"Kypros"
"Y_GE25","CY00",2005,4.3,"Kypros"
"Y_GE25","CZ",2005,6.8,"Czech Republic"
"Y_GE25","CZ0",2005,6.8,"Ceská republika"
"Y_GE25","CZ01",2005,3.1,"Praha"
"Y_GE25","CZ02",2005,4.6,"Strední Cechy"
"Y_GE25","CZ03",2005,4.3,"Jihozápad"
"Y_GE25","CZ04",2005,11.9,"Severozápad"
"Y_GE25","CZ05",2005,4.6,"Severovýchod"
"Y_GE25","CZ06",2005,6.5,"Jihovýchod"
"Y_GE25","CZ07",2005,8.5,"Strední Morava"
"Y_GE25","CZ08",2005,11.9,"Moravskoslezsko"
"Y_GE25","DE",2005,10.6,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2005,6.5,"Baden-Württemberg"
"Y_GE25","DE11",2005,6.8,"Stuttgart"
"Y_GE25","DE12",2005,7,"Karlsruhe"
"Y_GE25","DE13",2005,5.8,"Freiburg"
"Y_GE25","DE14",2005,6.2,"Tübingen"
"Y_GE25","DE2",2005,6.4,"Bayern"
"Y_GE25","DE21",2005,5.3,"Oberbayern"
"Y_GE25","DE22",2005,5.9,"Niederbayern"
"Y_GE25","DE23",2005,5.9,"Oberpfalz"
"Y_GE25","DE24",2005,9.3,"Oberfranken"
"Y_GE25","DE25",2005,8.1,"Mittelfranken"
"Y_GE25","DE26",2005,7,"Unterfranken"
"Y_GE25","DE27",2005,6.1,"Schwaben"
"Y_GE25","DE3",2005,18.8,"Berlin"
"Y_GE25","DE30",2005,18.8,"Berlin"
"Y_GE25","DE4",2005,17.6,"Brandenburg"
"Y_GE25","DE40",2005,17.6,"Brandenburg"
"Y_GE25","DE5",2005,16.3,"Bremen"
"Y_GE25","DE50",2005,16.3,"Bremen"
"Y_GE25","DE6",2005,10,"Hamburg"
"Y_GE25","DE60",2005,10,"Hamburg"
"Y_GE25","DE7",2005,8,"Hessen"
"Y_GE25","DE71",2005,7.7,"Darmstadt"
"Y_GE25","DE72",2005,8,"Gießen"
"Y_GE25","DE73",2005,8.9,"Kassel"
"Y_GE25","DE8",2005,21.4,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2005,21.4,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2005,9.8,"Niedersachsen"
"Y_GE25","DE91",2005,10.7,"Braunschweig"
"Y_GE25","DE92",2005,9.7,"Hannover"
"Y_GE25","DE93",2005,9,"Lüneburg"
"Y_GE25","DE94",2005,9.7,"Weser-Ems"
"Y_GE25","DEA",2005,9.8,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2005,10.1,"Düsseldorf"
"Y_GE25","DEA2",2005,8.8,"Köln"
"Y_GE25","DEA3",2005,8.8,"Münster"
"Y_GE25","DEA4",2005,9.5,"Detmold"
"Y_GE25","DEA5",2005,11.5,"Arnsberg"
"Y_GE25","DEB",2005,8.1,"Rheinland-Pfalz"
"Y_GE25","DEB1",2005,7.9,"Koblenz"
"Y_GE25","DEB2",2005,6.6,"Trier"
"Y_GE25","DEB3",2005,8.6,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2005,9.9,"Saarland"
"Y_GE25","DEC0",2005,9.9,"Saarland"
"Y_GE25","DED",2005,18.4,"Sachsen"
"Y_GE25","DED2",2005,18,"Dresden"
"Y_GE25","DED4",2005,18.2,"Chemnitz"
"Y_GE25","DED5",2005,19.6,"Leipzig"
"Y_GE25","DEE",2005,20,"Sachsen-Anhalt"
"Y_GE25","DEE0",2005,20,"Sachsen-Anhalt"
"Y_GE25","DEF",2005,9.7,"Schleswig-Holstein"
"Y_GE25","DEF0",2005,9.7,"Schleswig-Holstein"
"Y_GE25","DEG",2005,16.9,"Thüringen"
"Y_GE25","DEG0",2005,16.9,"Thüringen"
"Y_GE25","DK",2005,4.2,"Denmark"
"Y_GE25","DK0",2005,4.2,"Danmark"
"Y_GE25","EA17",2005,7.9,"Euro area (17 countries)"
"Y_GE25","EA18",2005,7.9,"Euro area (18 countries)"
"Y_GE25","EA19",2005,7.9,"Euro area (19 countries)"
"Y_GE25","EE",2005,7.2,"Estonia"
"Y_GE25","EE0",2005,7.2,"Eesti"
"Y_GE25","EE00",2005,7.2,"Eesti"
"Y_GE25","EL",2005,8.4,"Greece"
"Y_GE25","EL1",2005,9.8,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2005,9.6,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2005,9.5,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2005,15.5,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2005,8.5,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2005,8.4,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2005,9.6,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2005,7.1,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2005,9.3,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2005,8.5,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2005,7,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2005,7.6,"Attiki"
"Y_GE25","EL30",2005,7.6,"Attiki"
"Y_GE25","EL4",2005,7,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2005,7.3,"Voreio Aigaio"
"Y_GE25","EL42",2005,8.6,"Notio Aigaio"
"Y_GE25","EL43",2005,6.2,"Kriti"
"Y_GE25","ES",2005,7.7,"Spain"
"Y_GE25","ES1",2005,8.5,"Noroeste (ES)"
"Y_GE25","ES11",2005,8.6,"Galicia"
"Y_GE25","ES12",2005,8.6,"Principado de Asturias"
"Y_GE25","ES13",2005,7.4,"Cantabria"
"Y_GE25","ES2",2005,5.6,"Noreste (ES)"
"Y_GE25","ES21",2005,6.3,"País Vasco"
"Y_GE25","ES22",2005,4.7,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2005,5.3,"La Rioja"
"Y_GE25","ES24",2005,5,"Aragón"
"Y_GE25","ES3",2005,5.6,"Comunidad de Madrid"
"Y_GE25","ES30",2005,5.6,"Comunidad de Madrid"
"Y_GE25","ES4",2005,8.8,"Centro (ES)"
"Y_GE25","ES41",2005,7.5,"Castilla y León"
"Y_GE25","ES42",2005,7.8,"Castilla-la Mancha"
"Y_GE25","ES43",2005,13.7,"Extremadura"
"Y_GE25","ES5",2005,6.3,"Este (ES)"
"Y_GE25","ES51",2005,5.8,"Cataluña"
"Y_GE25","ES52",2005,7.4,"Comunidad Valenciana"
"Y_GE25","ES53",2005,5.6,"Illes Balears"
"Y_GE25","ES6",2005,11.2,"Sur (ES)"
"Y_GE25","ES61",2005,12,"Andalucía"
"Y_GE25","ES62",2005,6.8,"Región de Murcia"
"Y_GE25","ES63",2005,15.3,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2005,10.4,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2005,10,"Canarias (ES)"
"Y_GE25","ES70",2005,10,"Canarias (ES)"
"Y_GE25","EU15",2005,7,"European Union (15 countries)"
"Y_GE25","EU27",2005,7.6,"European Union (27 countries)"
"Y_GE25","EU28",2005,7.7,"European Union (28 countries)"
"Y_GE25","FI",2005,6.8,"Finland"
"Y_GE25","FI1",2005,6.8,"Manner-Suomi"
"Y_GE25","FI19",2005,7,"Länsi-Suomi"
"Y_GE25","FI1B",2005,4.8,"Helsinki-Uusimaa"
"Y_GE25","FI1C",2005,6.6,"Etelä-Suomi"
"Y_GE25","FI1D",2005,9.3,"Pohjois- ja Itä-Suomi"
"Y_GE25","FI2",2005,NA,"Åland"
"Y_GE25","FI20",2005,NA,"Åland"
"Y_GE25","FR",2005,7.5,"France"
"Y_GE25","FR1",2005,7.5,"Île de France"
"Y_GE25","FR10",2005,7.5,"Île de France"
"Y_GE25","FR2",2005,6.5,"Bassin Parisien"
"Y_GE25","FR21",2005,8.1,"Champagne-Ardenne"
"Y_GE25","FR22",2005,8.1,"Picardie"
"Y_GE25","FR23",2005,6.4,"Haute-Normandie"
"Y_GE25","FR24",2005,5.3,"Centre (FR)"
"Y_GE25","FR25",2005,6,"Basse-Normandie"
"Y_GE25","FR26",2005,5.6,"Bourgogne"
"Y_GE25","FR3",2005,10.2,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2005,10.2,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2005,6.5,"Est (FR)"
"Y_GE25","FR41",2005,7.9,"Lorraine"
"Y_GE25","FR42",2005,5.3,"Alsace"
"Y_GE25","FR43",2005,5.5,"Franche-Comté"
"Y_GE25","FR5",2005,5.9,"Ouest (FR)"
"Y_GE25","FR51",2005,5.7,"Pays de la Loire"
"Y_GE25","FR52",2005,5.7,"Bretagne"
"Y_GE25","FR53",2005,6.9,"Poitou-Charentes"
"Y_GE25","FR6",2005,6,"Sud-Ouest (FR)"
"Y_GE25","FR61",2005,6.3,"Aquitaine"
"Y_GE25","FR62",2005,5.9,"Midi-Pyrénées"
"Y_GE25","FR63",2005,4.7,"Limousin"
"Y_GE25","FR7",2005,6.6,"Centre-Est (FR)"
"Y_GE25","FR71",2005,6.7,"Rhône-Alpes"
"Y_GE25","FR72",2005,5.9,"Auvergne"
"Y_GE25","FR8",2005,9.1,"Méditerranée"
"Y_GE25","FR81",2005,10,"Languedoc-Roussillon"
"Y_GE25","FR82",2005,8.7,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2005,NA,"Corse"
"Y_GE25","FR9",2005,22.6,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2005,23.1,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2005,16.7,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2005,21.6,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2005,25.7,"Réunion (NUTS 2010)"
"Y_GE25","HR",2005,10.1,"Croatia"
"Y_GE25","HR0",2005,10.1,"Hrvatska"
"Y_GE25","HU",2005,6.1,"Hungary"
"Y_GE25","HU1",2005,4.4,"Közép-Magyarország"
"Y_GE25","HU10",2005,4.4,"Közép-Magyarország"
"Y_GE25","HU2",2005,6,"Dunántúl"
"Y_GE25","HU21",2005,5.6,"Közép-Dunántúl"
"Y_GE25","HU22",2005,5.2,"Nyugat-Dunántúl"
"Y_GE25","HU23",2005,7.3,"Dél-Dunántúl"
"Y_GE25","HU3",2005,7.7,"Alföld és Észak"
"Y_GE25","HU31",2005,8.8,"Észak-Magyarország"
"Y_GE25","HU32",2005,7.4,"Észak-Alföld"
"Y_GE25","HU33",2005,7,"Dél-Alföld"
"Y_GE25","IE",2005,3.5,"Ireland"
"Y_GE25","IE0",2005,3.5,"Éire/Ireland"
"Y_GE25","IE01",2005,3.5,"Border, Midland and Western"
"Y_GE25","IE02",2005,3.5,"Southern and Eastern"
"Y_GE25","IS",2005,1.6,"Iceland"
"Y_GE25","IS0",2005,1.6,"Ísland"
"Y_GE25","IS00",2005,1.6,"Ísland"
"Y_GE25","IT",2005,6.2,"Italy"
"Y_GE25","ITC",2005,3.6,"Nord-Ovest"
"Y_GE25","ITC1",2005,3.7,"Piemonte"
"Y_GE25","ITC2",2005,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2005,4.9,"Liguria"
"Y_GE25","ITC4",2005,3.3,"Lombardia"
"Y_GE25","ITF",2005,11.1,"Sud"
"Y_GE25","ITF1",2005,6.7,"Abruzzo"
"Y_GE25","ITF2",2005,8.1,"Molise"
"Y_GE25","ITF3",2005,12,"Campania"
"Y_GE25","ITF4",2005,11.9,"Puglia"
"Y_GE25","ITF5",2005,10.1,"Basilicata"
"Y_GE25","ITF6",2005,11.2,"Calabria"
"Y_GE25","ITG",2005,12.2,"Isole"
"Y_GE25","ITG1",2005,12.8,"Sicilia"
"Y_GE25","ITG2",2005,10.7,"Sardegna"
"Y_GE25","ITH",2005,3.4,"Nord-Est"
"Y_GE25","ITH1",2005,2.2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2005,3,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2005,3.5,"Veneto"
"Y_GE25","ITH4",2005,3.7,"Friuli-Venezia Giulia"
"Y_GE25","ITH5",2005,3.3,"Emilia-Romagna"
"Y_GE25","ITI",2005,5.3,"Centro (IT)"
"Y_GE25","ITI1",2005,4.6,"Toscana"
"Y_GE25","ITI2",2005,4.9,"Umbria"
"Y_GE25","ITI3",2005,4,"Marche"
"Y_GE25","ITI4",2005,6.3,"Lazio"
"Y_GE25","LT",2005,7.7,"Lithuania"
"Y_GE25","LT0",2005,7.7,"Lietuva"
"Y_GE25","LT00",2005,7.7,"Lietuva"
"Y_GE25","LU",2005,3.8,"Luxembourg"
"Y_GE25","LU0",2005,3.8,"Luxembourg"
"Y_GE25","LU00",2005,3.8,"Luxembourg"
"Y_GE25","LV",2005,9.3,"Latvia"
"Y_GE25","LV0",2005,9.3,"Latvija"
"Y_GE25","LV00",2005,9.3,"Latvija"
"Y_GE25","MT",2005,4.7,"Malta"
"Y_GE25","MT0",2005,4.7,"Malta"
"Y_GE25","MT00",2005,4.7,"Malta"
"Y_GE25","NL",2005,4.1,"Netherlands"
"Y_GE25","NL1",2005,4.9,"Noord-Nederland"
"Y_GE25","NL11",2005,6,"Groningen"
"Y_GE25","NL12",2005,3.9,"Friesland (NL)"
"Y_GE25","NL13",2005,4.9,"Drenthe"
"Y_GE25","NL2",2005,4.1,"Oost-Nederland"
"Y_GE25","NL21",2005,4.3,"Overijssel"
"Y_GE25","NL22",2005,3.7,"Gelderland"
"Y_GE25","NL23",2005,5.7,"Flevoland"
"Y_GE25","NL3",2005,4,"West-Nederland"
"Y_GE25","NL31",2005,3.2,"Utrecht"
"Y_GE25","NL32",2005,4.3,"Noord-Holland"
"Y_GE25","NL33",2005,4,"Zuid-Holland"
"Y_GE25","NL34",2005,2.8,"Zeeland"
"Y_GE25","NL4",2005,3.9,"Zuid-Nederland"
"Y_GE25","NL41",2005,3.4,"Noord-Brabant"
"Y_GE25","NL42",2005,4.9,"Limburg (NL)"
"Y_GE25","NO",2005,3.3,"Norway"
"Y_GE25","NO0",2005,3.3,"Norge"
"Y_GE25","NO01",2005,3.8,"Oslo og Akershus"
"Y_GE25","NO02",2005,3,"Hedmark og Oppland"
"Y_GE25","NO03",2005,3.5,"Sør-Østlandet"
"Y_GE25","NO04",2005,2.9,"Agder og Rogaland"
"Y_GE25","NO05",2005,3,"Vestlandet"
"Y_GE25","NO06",2005,2.5,"Trøndelag"
"Y_GE25","NO07",2005,3.5,"Nord-Norge"
"Y_GE25","PL",2005,15.1,"Poland"
"Y_GE25","PL1",2005,13.7,"Region Centralny"
"Y_GE25","PL11",2005,15.4,"Lódzkie"
"Y_GE25","PL12",2005,12.8,"Mazowieckie"
"Y_GE25","PL2",2005,14.6,"Region Poludniowy"
"Y_GE25","PL21",2005,12.4,"Malopolskie"
"Y_GE25","PL22",2005,16.1,"Slaskie"
"Y_GE25","PL3",2005,13.1,"Region Wschodni"
"Y_GE25","PL31",2005,12,"Lubelskie"
"Y_GE25","PL32",2005,13.2,"Podkarpackie"
"Y_GE25","PL33",2005,15.9,"Swietokrzyskie"
"Y_GE25","PL34",2005,12.2,"Podlaskie"
"Y_GE25","PL4",2005,16.1,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2005,13.9,"Wielkopolskie"
"Y_GE25","PL42",2005,20.1,"Zachodniopomorskie"
"Y_GE25","PL43",2005,16.8,"Lubuskie"
"Y_GE25","PL5",2005,18.7,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2005,20,"Dolnoslaskie"
"Y_GE25","PL52",2005,14.6,"Opolskie"
"Y_GE25","PL6",2005,16.8,"Region Pólnocny"
"Y_GE25","PL61",2005,16.6,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2005,18,"Warminsko-Mazurskie"
"Y_GE25","PL63",2005,16.1,"Pomorskie"
"Y_GE25","PT",2005,6.6,"Portugal"
"Y_GE25","PT1",2005,6.8,"Continente"
"Y_GE25","PT11",2005,7.8,"Norte"
"Y_GE25","PT15",2005,5.4,"Algarve"
"Y_GE25","PT16",2005,4.2,"Centro (PT)"
"Y_GE25","PT17",2005,7.7,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2005,7.8,"Alentejo"
"Y_GE25","PT2",2005,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2005,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2005,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2005,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2005,5.6,"Romania"
"Y_GE25","RO1",2005,5.6,"Macroregiunea unu"
"Y_GE25","RO11",2005,4.3,"Nord-Vest"
"Y_GE25","RO12",2005,7,"Centru"
"Y_GE25","RO2",2005,5.1,"Macroregiunea doi"
"Y_GE25","RO21",2005,4.2,"Nord-Est"
"Y_GE25","RO22",2005,6.3,"Sud-Est"
"Y_GE25","RO3",2005,6.5,"Macroregiunea trei"
"Y_GE25","RO31",2005,7.3,"Sud - Muntenia"
"Y_GE25","RO32",2005,5.4,"Bucuresti - Ilfov"
"Y_GE25","RO4",2005,5.4,"Macroregiunea patru"
"Y_GE25","RO41",2005,5.3,"Sud-Vest Oltenia"
"Y_GE25","RO42",2005,5.4,"Vest"
"Y_GE25","SE",2005,5.8,"Sweden"
"Y_GE25","SE1",2005,5.6,"Östra Sverige"
"Y_GE25","SE11",2005,5.2,"Stockholm"
"Y_GE25","SE12",2005,6.2,"Östra Mellansverige"
"Y_GE25","SE2",2005,5.6,"Södra Sverige"
"Y_GE25","SE21",2005,4.3,"Småland med öarna"
"Y_GE25","SE22",2005,7,"Sydsverige"
"Y_GE25","SE23",2005,5.1,"Västsverige"
"Y_GE25","SE3",2005,6.7,"Norra Sverige"
"Y_GE25","SE31",2005,6.9,"Norra Mellansverige"
"Y_GE25","SE32",2005,6.8,"Mellersta Norrland"
"Y_GE25","SE33",2005,6.5,"Övre Norrland"
"Y_GE25","SI",2005,5.4,"Slovenia"
"Y_GE25","SI0",2005,5.4,"Slovenija"
"Y_GE25","SI01",2005,6.3,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2005,4.4,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2005,14.4,"Slovakia"
"Y_GE25","SK0",2005,14.4,"Slovensko"
"Y_GE25","SK01",2005,4.8,"Bratislavský kraj"
"Y_GE25","SK02",2005,11.2,"Západné Slovensko"
"Y_GE25","SK03",2005,17.4,"Stredné Slovensko"
"Y_GE25","SK04",2005,20.2,"Východné Slovensko"
"Y_GE25","UK",2005,3.3,"United Kingdom"
"Y_GE25","UKC",2005,4,"North East (UK)"
"Y_GE25","UKC1",2005,4,"Tees Valley and Durham"
"Y_GE25","UKC2",2005,4.1,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2005,3,"North West (UK)"
"Y_GE25","UKD1",2005,2,"Cumbria"
"Y_GE25","UKD3",2005,3.3,"Greater Manchester"
"Y_GE25","UKD4",2005,2.8,"Lancashire"
"Y_GE25","UKD6",2005,2.4,"Cheshire"
"Y_GE25","UKD7",2005,3.6,"Merseyside"
"Y_GE25","UKE",2005,3,"Yorkshire and The Humber"
"Y_GE25","UKE1",2005,3.7,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2005,2,"North Yorkshire"
"Y_GE25","UKE3",2005,3.6,"South Yorkshire"
"Y_GE25","UKE4",2005,2.7,"West Yorkshire"
"Y_GE25","UKF",2005,3,"East Midlands (UK)"
"Y_GE25","UKF1",2005,3.1,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2005,3.1,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2005,2.6,"Lincolnshire"
"Y_GE25","UKG",2005,3.3,"West Midlands (UK)"
"Y_GE25","UKG1",2005,1.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2005,2.7,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2005,4.4,"West Midlands"
"Y_GE25","UKH",2005,2.8,"East of England"
"Y_GE25","UKH1",2005,3,"East Anglia"
"Y_GE25","UKH2",2005,2.7,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2005,2.6,"Essex"
"Y_GE25","UKI",2005,5.1,"London"
"Y_GE25","UKI1",2005,5.9,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2005,4.6,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2005,2.7,"South East (UK)"
"Y_GE25","UKJ1",2005,2.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2005,2.9,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2005,2.5,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2005,3.1,"Kent"
"Y_GE25","UKK",2005,2.4,"South West (UK)"
"Y_GE25","UKK1",2005,2.2,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2005,2.9,"Dorset and Somerset"
"Y_GE25","UKK3",2005,2.3,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2005,2.5,"Devon"
"Y_GE25","UKL",2005,2.9,"Wales"
"Y_GE25","UKL1",2005,3.2,"West Wales and The Valleys"
"Y_GE25","UKL2",2005,2.4,"East Wales"
"Y_GE25","UKM",2005,3.8,"Scotland"
"Y_GE25","UKM2",2005,3.5,"Eastern Scotland"
"Y_GE25","UKM3",2005,4.6,"South Western Scotland"
"Y_GE25","UKM5",2005,2.5,"North Eastern Scotland"
"Y_GE25","UKM6",2005,2.6,"Highlands and Islands"
"Y_GE25","UKN",2005,3.4,"Northern Ireland (UK)"
"Y_GE25","UKN0",2005,3.4,"Northern Ireland (UK)"
"Y15-24","AT",2004,12.1,"Austria"
"Y15-24","AT1",2004,16.8,"Ostösterreich"
"Y15-24","AT11",2004,NA,"Burgenland (AT)"
"Y15-24","AT12",2004,12.3,"Niederösterreich"
"Y15-24","AT13",2004,22.1,"Wien"
"Y15-24","AT2",2004,8.4,"Südösterreich"
"Y15-24","AT21",2004,NA,"Kärnten"
"Y15-24","AT22",2004,7.5,"Steiermark"
"Y15-24","AT3",2004,9.7,"Westösterreich"
"Y15-24","AT31",2004,11.5,"Oberösterreich"
"Y15-24","AT32",2004,NA,"Salzburg"
"Y15-24","AT33",2004,NA,"Tirol"
"Y15-24","AT34",2004,NA,"Vorarlberg"
"Y15-24","BE",2004,17.5,"Belgium"
"Y15-24","BE1",2004,19.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2004,19.2,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2004,11.9,"Vlaams Gewest"
"Y15-24","BE21",2004,14.5,"Prov. Antwerpen"
"Y15-24","BE22",2004,14.4,"Prov. Limburg (BE)"
"Y15-24","BE23",2004,13,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2004,NA,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2004,NA,"Prov. West-Vlaanderen"
"Y15-24","BE3",2004,28.9,"Région wallonne"
"Y15-24","BE31",2004,NA,"Prov. Brabant Wallon"
"Y15-24","BE32",2004,35,"Prov. Hainaut"
"Y15-24","BE33",2004,27.2,"Prov. Liège"
"Y15-24","BE34",2004,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2004,NA,"Prov. Namur"
"Y15-24","BG",2004,24.5,"Bulgaria"
"Y15-24","BG3",2004,29.5,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2004,24.5,"Severozapaden"
"Y15-24","BG32",2004,31.6,"Severen tsentralen"
"Y15-24","BG33",2004,32.9,"Severoiztochen"
"Y15-24","BG34",2004,27.4,"Yugoiztochen"
"Y15-24","BG4",2004,19.6,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2004,17.7,"Yugozapaden"
"Y15-24","BG42",2004,22.4,"Yuzhen tsentralen"
"Y15-24","CH",2004,7.7,"Switzerland"
"Y15-24","CH0",2004,7.7,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2004,10.2,"Région lémanique"
"Y15-24","CH02",2004,6.6,"Espace Mittelland"
"Y15-24","CH03",2004,7.2,"Nordwestschweiz"
"Y15-24","CH04",2004,11.5,"Zürich"
"Y15-24","CH05",2004,5.6,"Ostschweiz"
"Y15-24","CH06",2004,4,"Zentralschweiz"
"Y15-24","CH07",2004,NA,"Ticino"
"Y15-24","CY",2004,8.7,"Cyprus"
"Y15-24","CY0",2004,8.7,"Kypros"
"Y15-24","CY00",2004,8.7,"Kypros"
"Y15-24","CZ",2004,19.9,"Czech Republic"
"Y15-24","CZ0",2004,19.9,"Ceská republika"
"Y15-24","CZ01",2004,9.1,"Praha"
"Y15-24","CZ02",2004,9.6,"Strední Cechy"
"Y15-24","CZ03",2004,11.5,"Jihozápad"
"Y15-24","CZ04",2004,26.3,"Severozápad"
"Y15-24","CZ05",2004,16.6,"Severovýchod"
"Y15-24","CZ06",2004,20.4,"Jihovýchod"
"Y15-24","CZ07",2004,27,"Strední Morava"
"Y15-24","CZ08",2004,33.3,"Moravskoslezsko"
"Y15-24","DE",2004,13,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2004,9.6,"Baden-Württemberg"
"Y15-24","DE11",2004,8.6,"Stuttgart"
"Y15-24","DE12",2004,9.4,"Karlsruhe"
"Y15-24","DE13",2004,11.2,"Freiburg"
"Y15-24","DE14",2004,9.9,"Tübingen"
"Y15-24","DE2",2004,8.9,"Bayern"
"Y15-24","DE21",2004,7.7,"Oberbayern"
"Y15-24","DE22",2004,8.5,"Niederbayern"
"Y15-24","DE23",2004,NA,"Oberpfalz"
"Y15-24","DE24",2004,13.4,"Oberfranken"
"Y15-24","DE25",2004,7.9,"Mittelfranken"
"Y15-24","DE26",2004,12.5,"Unterfranken"
"Y15-24","DE27",2004,8.2,"Schwaben"
"Y15-24","DE3",2004,21,"Berlin"
"Y15-24","DE30",2004,21,"Berlin"
"Y15-24","DE4",2004,22.6,"Brandenburg"
"Y15-24","DE40",2004,22.6,"Brandenburg"
"Y15-24","DE5",2004,20.1,"Bremen"
"Y15-24","DE50",2004,20.1,"Bremen"
"Y15-24","DE6",2004,14.3,"Hamburg"
"Y15-24","DE60",2004,14.3,"Hamburg"
"Y15-24","DE7",2004,12.2,"Hessen"
"Y15-24","DE71",2004,12.2,"Darmstadt"
"Y15-24","DE72",2004,12.7,"Gießen"
"Y15-24","DE73",2004,11.7,"Kassel"
"Y15-24","DE8",2004,19.2,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2004,19.2,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2004,11.7,"Niedersachsen"
"Y15-24","DE91",2004,10.6,"Braunschweig"
"Y15-24","DE92",2004,13.8,"Hannover"
"Y15-24","DE93",2004,12.8,"Lüneburg"
"Y15-24","DE94",2004,10,"Weser-Ems"
"Y15-24","DEA",2004,12.2,"Nordrhein-Westfalen"
"Y15-24","DEA1",2004,12.5,"Düsseldorf"
"Y15-24","DEA2",2004,9.4,"Köln"
"Y15-24","DEA3",2004,13.1,"Münster"
"Y15-24","DEA4",2004,14,"Detmold"
"Y15-24","DEA5",2004,12.9,"Arnsberg"
"Y15-24","DEB",2004,12.4,"Rheinland-Pfalz"
"Y15-24","DEB1",2004,13.3,"Koblenz"
"Y15-24","DEB2",2004,NA,"Trier"
"Y15-24","DEB3",2004,11.6,"Rheinhessen-Pfalz"
"Y15-24","DEC",2004,12.7,"Saarland"
"Y15-24","DEC0",2004,12.7,"Saarland"
"Y15-24","DED",2004,17.1,"Sachsen"
"Y15-24","DED2",2004,18,"Dresden"
"Y15-24","DEE",2004,17.7,"Sachsen-Anhalt"
"Y15-24","DEE0",2004,17.7,"Sachsen-Anhalt"
"Y15-24","DEF",2004,14.8,"Schleswig-Holstein"
"Y15-24","DEF0",2004,14.8,"Schleswig-Holstein"
"Y15-24","DEG",2004,14.1,"Thüringen"
"Y15-24","DEG0",2004,14.1,"Thüringen"
"Y15-24","DK",2004,7.8,"Denmark"
"Y15-24","DK0",2004,7.8,"Danmark"
"Y15-24","EA17",2004,18,"Euro area (17 countries)"
"Y15-24","EA18",2004,18.1,"Euro area (18 countries)"
"Y15-24","EA19",2004,18.1,"Euro area (19 countries)"
"Y15-24","EE",2004,25.7,"Estonia"
"Y15-24","EE0",2004,25.7,"Eesti"
"Y15-24","EE00",2004,25.7,"Eesti"
"Y15-24","EL",2004,26.1,"Greece"
"Y15-24","EL1",2004,32,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2004,31,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2004,31.9,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2004,52.8,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2004,25.7,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2004,29.8,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2004,34,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2004,23.8,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2004,28.2,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2004,30.8,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2004,30.8,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2004,21.9,"Attiki"
"Y15-24","EL30",2004,21.9,"Attiki"
"Y15-24","EL4",2004,19.1,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2004,21.8,"Voreio Aigaio"
"Y15-24","EL42",2004,20.3,"Notio Aigaio"
"Y15-24","EL43",2004,17.6,"Kriti"
"Y15-24","ES",2004,22.5,"Spain"
"Y15-24","ES1",2004,27.6,"Noroeste (ES)"
"Y15-24","ES11",2004,27.8,"Galicia"
"Y15-24","ES12",2004,30.1,"Principado de Asturias"
"Y15-24","ES13",2004,22.4,"Cantabria"
"Y15-24","ES2",2004,18.6,"Noreste (ES)"
"Y15-24","ES21",2004,24.8,"País Vasco"
"Y15-24","ES22",2004,12.7,"Comunidad Foral de Navarra"
"Y15-24","ES23",2004,NA,"La Rioja"
"Y15-24","ES24",2004,13.8,"Aragón"
"Y15-24","ES3",2004,13.8,"Comunidad de Madrid"
"Y15-24","ES30",2004,13.8,"Comunidad de Madrid"
"Y15-24","ES4",2004,21.1,"Centro (ES)"
"Y15-24","ES41",2004,22.8,"Castilla y León"
"Y15-24","ES42",2004,15.3,"Castilla-la Mancha"
"Y15-24","ES43",2004,28.8,"Extremadura"
"Y15-24","ES5",2004,21.3,"Este (ES)"
"Y15-24","ES51",2004,23,"Cataluña"
"Y15-24","ES52",2004,19.7,"Comunidad Valenciana"
"Y15-24","ES53",2004,17.4,"Illes Balears"
"Y15-24","ES6",2004,27.7,"Sur (ES)"
"Y15-24","ES61",2004,28.8,"Andalucía"
"Y15-24","ES62",2004,21.2,"Región de Murcia"
"Y15-24","ES63",2004,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2004,NA,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2004,28.2,"Canarias (ES)"
"Y15-24","ES70",2004,28.2,"Canarias (ES)"
"Y15-24","EU15",2004,16.1,"European Union (15 countries)"
"Y15-24","EU27",2004,18.7,"European Union (27 countries)"
"Y15-24","EU28",2004,18.8,"European Union (28 countries)"
"Y15-24","FI",2004,27.5,"Finland"
"Y15-24","FI1",2004,27.6,"Manner-Suomi"
"Y15-24","FI19",2004,27.2,"Länsi-Suomi"
"Y15-24","FI2",2004,NA,"Åland"
"Y15-24","FI20",2004,NA,"Åland"
"Y15-24","FR",2004,20.7,"France"
"Y15-24","FR1",2004,18.7,"Île de France"
"Y15-24","FR10",2004,18.7,"Île de France"
"Y15-24","FR2",2004,21.3,"Bassin Parisien"
"Y15-24","FR21",2004,NA,"Champagne-Ardenne"
"Y15-24","FR22",2004,NA,"Picardie"
"Y15-24","FR23",2004,NA,"Haute-Normandie"
"Y15-24","FR24",2004,NA,"Centre (FR)"
"Y15-24","FR25",2004,NA,"Basse-Normandie"
"Y15-24","FR26",2004,NA,"Bourgogne"
"Y15-24","FR3",2004,28.9,"Nord - Pas-de-Calais"
"Y15-24","FR30",2004,28.9,"Nord - Pas-de-Calais"
"Y15-24","FR4",2004,22.7,"Est (FR)"
"Y15-24","FR41",2004,NA,"Lorraine"
"Y15-24","FR42",2004,NA,"Alsace"
"Y15-24","FR43",2004,NA,"Franche-Comté"
"Y15-24","FR5",2004,15.4,"Ouest (FR)"
"Y15-24","FR51",2004,NA,"Pays de la Loire"
"Y15-24","FR52",2004,NA,"Bretagne"
"Y15-24","FR53",2004,NA,"Poitou-Charentes"
"Y15-24","FR6",2004,20,"Sud-Ouest (FR)"
"Y15-24","FR61",2004,NA,"Aquitaine"
"Y15-24","FR62",2004,NA,"Midi-Pyrénées"
"Y15-24","FR63",2004,NA,"Limousin"
"Y15-24","FR7",2004,15.1,"Centre-Est (FR)"
"Y15-24","FR71",2004,14.2,"Rhône-Alpes"
"Y15-24","FR72",2004,NA,"Auvergne"
"Y15-24","FR8",2004,20.5,"Méditerranée"
"Y15-24","FR81",2004,NA,"Languedoc-Roussillon"
"Y15-24","FR82",2004,18.3,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2004,NA,"Corse"
"Y15-24","FR9",2004,54.8,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2004,55.9,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2004,49.3,"Martinique (NUTS 2010)"
"Y15-24","FR93",2004,49.3,"Guyane (NUTS 2010)"
"Y15-24","FR94",2004,56.6,"Réunion (NUTS 2010)"
"Y15-24","HR",2004,32.8,"Croatia"
"Y15-24","HR0",2004,32.8,"Hrvatska"
"Y15-24","HU",2004,14.4,"Hungary"
"Y15-24","HU1",2004,11.9,"Közép-Magyarország"
"Y15-24","HU10",2004,11.9,"Közép-Magyarország"
"Y15-24","HU2",2004,12.7,"Dunántúl"
"Y15-24","HU21",2004,12.2,"Közép-Dunántúl"
"Y15-24","HU22",2004,9.3,"Nyugat-Dunántúl"
"Y15-24","HU23",2004,17.4,"Dél-Dunántúl"
"Y15-24","HU3",2004,17.7,"Alföld és Észak"
"Y15-24","HU31",2004,20.7,"Észak-Magyarország"
"Y15-24","HU32",2004,16.2,"Észak-Alföld"
"Y15-24","HU33",2004,16.5,"Dél-Alföld"
"Y15-24","IE",2004,8.3,"Ireland"
"Y15-24","IE0",2004,8.3,"Éire/Ireland"
"Y15-24","IE01",2004,8.6,"Border, Midland and Western"
"Y15-24","IE02",2004,8.2,"Southern and Eastern"
"Y15-24","IS",2004,12.1,"Iceland"
"Y15-24","IS0",2004,12.1,"Ísland"
"Y15-24","IS00",2004,12.1,"Ísland"
"Y15-24","IT",2004,24.4,"Italy"
"Y15-24","ITC",2004,13.2,"Nord-Ovest"
"Y15-24","ITC1",2004,15,"Piemonte"
"Y15-24","ITC2",2004,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2004,19.6,"Liguria"
"Y15-24","ITC4",2004,11.9,"Lombardia"
"Y15-24","ITF",2004,37.9,"Sud"
"Y15-24","ITF1",2004,29,"Abruzzo"
"Y15-24","ITF2",2004,35,"Molise"
"Y15-24","ITF3",2004,39.7,"Campania"
"Y15-24","ITF4",2004,34.9,"Puglia"
"Y15-24","ITF5",2004,32.5,"Basilicata"
"Y15-24","ITF6",2004,46.3,"Calabria"
"Y15-24","ITG",2004,40.9,"Isole"
"Y15-24","ITG1",2004,42.1,"Sicilia"
"Y15-24","ITG2",2004,37.9,"Sardegna"
"Y15-24","ITH",2004,12.9,"Nord-Est"
"Y15-24","ITH1",2004,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2004,NA,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2004,11.7,"Veneto"
"Y15-24","ITH4",2004,14.2,"Friuli-Venezia Giulia"
"Y15-24","ITI",2004,23.1,"Centro (IT)"
"Y15-24","ITI1",2004,18.2,"Toscana"
"Y15-24","ITI2",2004,16.1,"Umbria"
"Y15-24","ITI4",2004,30.5,"Lazio"
"Y15-24","LT",2004,20.3,"Lithuania"
"Y15-24","LT0",2004,20.3,"Lietuva"
"Y15-24","LT00",2004,20.3,"Lietuva"
"Y15-24","LU",2004,16.9,"Luxembourg"
"Y15-24","LU0",2004,16.9,"Luxembourg"
"Y15-24","LU00",2004,16.9,"Luxembourg"
"Y15-24","LV",2004,21.8,"Latvia"
"Y15-24","LV0",2004,21.8,"Latvija"
"Y15-24","LV00",2004,21.8,"Latvija"
"Y15-24","MT",2004,18.3,"Malta"
"Y15-24","MT0",2004,18.3,"Malta"
"Y15-24","MT00",2004,18.3,"Malta"
"Y15-24","NL",2004,8,"Netherlands"
"Y15-24","NL1",2004,8.6,"Noord-Nederland"
"Y15-24","NL11",2004,8.6,"Groningen"
"Y15-24","NL12",2004,7.7,"Friesland (NL)"
"Y15-24","NL13",2004,9.8,"Drenthe"
"Y15-24","NL2",2004,8.8,"Oost-Nederland"
"Y15-24","NL21",2004,9,"Overijssel"
"Y15-24","NL22",2004,7.2,"Gelderland"
"Y15-24","NL23",2004,16,"Flevoland"
"Y15-24","NL3",2004,8,"West-Nederland"
"Y15-24","NL31",2004,7.1,"Utrecht"
"Y15-24","NL32",2004,10,"Noord-Holland"
"Y15-24","NL33",2004,7.3,"Zuid-Holland"
"Y15-24","NL34",2004,4.9,"Zeeland"
"Y15-24","NL4",2004,6.9,"Zuid-Nederland"
"Y15-24","NL41",2004,6.8,"Noord-Brabant"
"Y15-24","NL42",2004,7.4,"Limburg (NL)"
"Y15-24","NO",2004,12.8,"Norway"
"Y15-24","NO0",2004,12.8,"Norge"
"Y15-24","NO01",2004,11.8,"Oslo og Akershus"
"Y15-24","NO02",2004,14.3,"Hedmark og Oppland"
"Y15-24","NO03",2004,13,"Sør-Østlandet"
"Y15-24","NO04",2004,13.1,"Agder og Rogaland"
"Y15-24","NO05",2004,11.4,"Vestlandet"
"Y15-24","NO06",2004,10.4,"Trøndelag"
"Y15-24","NO07",2004,16.9,"Nord-Norge"
"Y15-24","PL",2004,40.1,"Poland"
"Y15-24","PL1",2004,36.1,"Region Centralny"
"Y15-24","PL11",2004,38.5,"Lódzkie"
"Y15-24","PL12",2004,34.6,"Mazowieckie"
"Y15-24","PL2",2004,43,"Region Poludniowy"
"Y15-24","PL21",2004,41.4,"Malopolskie"
"Y15-24","PL22",2004,44.1,"Slaskie"
"Y15-24","PL3",2004,36.7,"Region Wschodni"
"Y15-24","PL31",2004,37.5,"Lubelskie"
"Y15-24","PL32",2004,35.4,"Podkarpackie"
"Y15-24","PL33",2004,39.8,"Swietokrzyskie"
"Y15-24","PL34",2004,33.5,"Podlaskie"
"Y15-24","PL4",2004,39.8,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2004,36.4,"Wielkopolskie"
"Y15-24","PL42",2004,39.1,"Zachodniopomorskie"
"Y15-24","PL43",2004,52.5,"Lubuskie"
"Y15-24","PL5",2004,47.5,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2004,48.7,"Dolnoslaskie"
"Y15-24","PL52",2004,42.5,"Opolskie"
"Y15-24","PL6",2004,40.2,"Region Pólnocny"
"Y15-24","PL61",2004,39.9,"Kujawsko-Pomorskie"
"Y15-24","PL62",2004,47.4,"Warminsko-Mazurskie"
"Y15-24","PL63",2004,36.2,"Pomorskie"
"Y15-24","PT",2004,14.1,"Portugal"
"Y15-24","PT1",2004,14.4,"Continente"
"Y15-24","PT11",2004,14.2,"Norte"
"Y15-24","PT15",2004,NA,"Algarve"
"Y15-24","PT16",2004,8.7,"Centro (PT)"
"Y15-24","PT17",2004,17.6,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2004,23.4,"Alentejo"
"Y15-24","PT2",2004,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2004,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2004,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2004,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2004,22.3,"Romania"
"Y15-24","RO1",2004,21.4,"Macroregiunea unu"
"Y15-24","RO11",2004,19,"Nord-Vest"
"Y15-24","RO12",2004,24.1,"Centru"
"Y15-24","RO2",2004,19.2,"Macroregiunea doi"
"Y15-24","RO21",2004,17.6,"Nord-Est"
"Y15-24","RO22",2004,21.7,"Sud-Est"
"Y15-24","RO3",2004,28.3,"Macroregiunea trei"
"Y15-24","RO31",2004,29,"Sud - Muntenia"
"Y15-24","RO32",2004,27.2,"Bucuresti - Ilfov"
"Y15-24","RO4",2004,21,"Macroregiunea patru"
"Y15-24","RO41",2004,16.8,"Sud-Vest Oltenia"
"Y15-24","RO42",2004,25.4,"Vest"
"Y15-24","SE",2004,18.5,"Sweden"
"Y15-24","SE1",2004,18.8,"Östra Sverige"
"Y15-24","SE11",2004,17.6,"Stockholm"
"Y15-24","SE12",2004,20.2,"Östra Mellansverige"
"Y15-24","SE2",2004,17.6,"Södra Sverige"
"Y15-24","SE21",2004,15.9,"Småland med öarna"
"Y15-24","SE22",2004,20.7,"Sydsverige"
"Y15-24","SE23",2004,16.3,"Västsverige"
"Y15-24","SE3",2004,20.4,"Norra Sverige"
"Y15-24","SE31",2004,21,"Norra Mellansverige"
"Y15-24","SE32",2004,22.3,"Mellersta Norrland"
"Y15-24","SE33",2004,18.3,"Övre Norrland"
"Y15-24","SI",2004,14,"Slovenia"
"Y15-24","SI0",2004,14,"Slovenija"
"Y15-24","SI01",2004,16.6,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2004,10.6,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2004,32.8,"Slovakia"
"Y15-24","SK0",2004,32.8,"Slovensko"
"Y15-24","SK01",2004,19.7,"Bratislavský kraj"
"Y15-24","SK02",2004,24.6,"Západné Slovensko"
"Y15-24","SK03",2004,37.7,"Stredné Slovensko"
"Y15-24","SK04",2004,42.8,"Východné Slovensko"
"Y15-24","UK",2004,10.7,"United Kingdom"
"Y15-24","UKC",2004,12.9,"North East (UK)"
"Y15-24","UKC1",2004,13.8,"Tees Valley and Durham"
"Y15-24","UKC2",2004,12.1,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2004,11.1,"North West (UK)"
"Y15-24","UKD1",2004,NA,"Cumbria"
"Y15-24","UKD3",2004,13,"Greater Manchester"
"Y15-24","UKD4",2004,10.1,"Lancashire"
"Y15-24","UKE",2004,9.3,"Yorkshire and The Humber"
"Y15-24","UKE1",2004,NA,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2004,NA,"North Yorkshire"
"Y15-24","UKE3",2004,NA,"South Yorkshire"
"Y15-24","UKE4",2004,9.9,"West Yorkshire"
"Y15-24","UKF",2004,7.5,"East Midlands (UK)"
"Y15-24","UKF1",2004,6.9,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2004,8.4,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2004,NA,"Lincolnshire"
"Y15-24","UKG",2004,12.2,"West Midlands (UK)"
"Y15-24","UKG1",2004,NA,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2004,9.1,"Shropshire and Staffordshire"
"Y15-24","UKG3",2004,15.6,"West Midlands"
"Y15-24","UKH",2004,10,"East of England"
"Y15-24","UKH1",2004,11.6,"East Anglia"
"Y15-24","UKH2",2004,8.7,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2004,9.6,"Essex"
"Y15-24","UKI",2004,15.3,"London"
"Y15-24","UKI1",2004,19.8,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2004,12.2,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2004,8.4,"South East (UK)"
"Y15-24","UKJ1",2004,9.4,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2004,7,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2004,8.1,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2004,9.3,"Kent"
"Y15-24","UKK",2004,7.8,"South West (UK)"
"Y15-24","UKK1",2004,8.1,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2004,NA,"Dorset and Somerset"
"Y15-24","UKK3",2004,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2004,NA,"Devon"
"Y15-24","UKL",2004,10.4,"Wales"
"Y15-24","UKL1",2004,13.3,"West Wales and The Valleys"
"Y15-24","UKL2",2004,NA,"East Wales"
"Y15-24","UKM",2004,13,"Scotland"
"Y15-24","UKM2",2004,12.2,"Eastern Scotland"
"Y15-24","UKM3",2004,14.7,"South Western Scotland"
"Y15-24","UKM5",2004,NA,"North Eastern Scotland"
"Y15-24","UKM6",2004,NA,"Highlands and Islands"
"Y15-24","UKN",2004,9.8,"Northern Ireland (UK)"
"Y15-24","UKN0",2004,9.8,"Northern Ireland (UK)"
"Y20-64","AT",2004,5.4,"Austria"
"Y20-64","AT1",2004,6.9,"Ostösterreich"
"Y20-64","AT11",2004,5,"Burgenland (AT)"
"Y20-64","AT12",2004,4.1,"Niederösterreich"
"Y20-64","AT13",2004,9.8,"Wien"
"Y20-64","AT2",2004,5,"Südösterreich"
"Y20-64","AT21",2004,6,"Kärnten"
"Y20-64","AT22",2004,4.5,"Steiermark"
"Y20-64","AT3",2004,4,"Westösterreich"
"Y20-64","AT31",2004,4.5,"Oberösterreich"
"Y20-64","AT32",2004,4.2,"Salzburg"
"Y20-64","AT33",2004,2.6,"Tirol"
"Y20-64","AT34",2004,3.9,"Vorarlberg"
"Y20-64","BE",2004,7.1,"Belgium"
"Y20-64","BE1",2004,13.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2004,13.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2004,4.4,"Vlaams Gewest"
"Y20-64","BE21",2004,5.2,"Prov. Antwerpen"
"Y20-64","BE22",2004,5.6,"Prov. Limburg (BE)"
"Y20-64","BE23",2004,4,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2004,4,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2004,3,"Prov. West-Vlaanderen"
"Y20-64","BE3",2004,10.6,"Région wallonne"
"Y20-64","BE31",2004,6.3,"Prov. Brabant Wallon"
"Y20-64","BE32",2004,12.2,"Prov. Hainaut"
"Y20-64","BE33",2004,12.9,"Prov. Liège"
"Y20-64","BE34",2004,6.7,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2004,7.5,"Prov. Namur"
"Y20-64","BG",2004,11.8,"Bulgaria"
"Y20-64","BG3",2004,14.3,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2004,12.3,"Severozapaden"
"Y20-64","BG32",2004,14.7,"Severen tsentralen"
"Y20-64","BG33",2004,17.6,"Severoiztochen"
"Y20-64","BG34",2004,12.6,"Yugoiztochen"
"Y20-64","BG4",2004,9.2,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2004,9,"Yugozapaden"
"Y20-64","BG42",2004,9.5,"Yuzhen tsentralen"
"Y20-64","CH",2004,4.2,"Switzerland"
"Y20-64","CH0",2004,4.2,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2004,5.6,"Région lémanique"
"Y20-64","CH02",2004,3.6,"Espace Mittelland"
"Y20-64","CH03",2004,3.7,"Nordwestschweiz"
"Y20-64","CH04",2004,4.8,"Zürich"
"Y20-64","CH05",2004,3.5,"Ostschweiz"
"Y20-64","CH06",2004,3.4,"Zentralschweiz"
"Y20-64","CH07",2004,5.5,"Ticino"
"Y20-64","CY",2004,4.3,"Cyprus"
"Y20-64","CY0",2004,4.3,"Kypros"
"Y20-64","CY00",2004,4.3,"Kypros"
"Y20-64","CZ",2004,8,"Czech Republic"
"Y20-64","CZ0",2004,8,"Ceská republika"
"Y20-64","CZ01",2004,3.9,"Praha"
"Y20-64","CZ02",2004,5.4,"Strední Cechy"
"Y20-64","CZ03",2004,5.7,"Jihozápad"
"Y20-64","CZ04",2004,11.5,"Severozápad"
"Y20-64","CZ05",2004,6.4,"Severovýchod"
"Y20-64","CZ06",2004,7.7,"Jihovýchod"
"Y20-64","CZ07",2004,9.7,"Strední Morava"
"Y20-64","CZ08",2004,14.2,"Moravskoslezsko"
"Y20-64","DE",2004,10.9,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2004,6.6,"Baden-Württemberg"
"Y20-64","DE11",2004,6.8,"Stuttgart"
"Y20-64","DE12",2004,6.9,"Karlsruhe"
"Y20-64","DE13",2004,6.4,"Freiburg"
"Y20-64","DE14",2004,6.2,"Tübingen"
"Y20-64","DE2",2004,6.9,"Bayern"
"Y20-64","DE21",2004,5.3,"Oberbayern"
"Y20-64","DE22",2004,6.4,"Niederbayern"
"Y20-64","DE23",2004,7.2,"Oberpfalz"
"Y20-64","DE24",2004,10,"Oberfranken"
"Y20-64","DE25",2004,8.8,"Mittelfranken"
"Y20-64","DE26",2004,7.5,"Unterfranken"
"Y20-64","DE27",2004,6.9,"Schwaben"
"Y20-64","DE3",2004,19.2,"Berlin"
"Y20-64","DE30",2004,19.2,"Berlin"
"Y20-64","DE4",2004,19.6,"Brandenburg"
"Y20-64","DE40",2004,19.6,"Brandenburg"
"Y20-64","DE5",2004,14.8,"Bremen"
"Y20-64","DE50",2004,14.8,"Bremen"
"Y20-64","DE6",2004,10.7,"Hamburg"
"Y20-64","DE60",2004,10.7,"Hamburg"
"Y20-64","DE7",2004,7.9,"Hessen"
"Y20-64","DE71",2004,7.8,"Darmstadt"
"Y20-64","DE72",2004,8.6,"Gießen"
"Y20-64","DE73",2004,7.7,"Kassel"
"Y20-64","DE8",2004,23,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2004,23,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2004,9.6,"Niedersachsen"
"Y20-64","DE91",2004,10.6,"Braunschweig"
"Y20-64","DE92",2004,10,"Hannover"
"Y20-64","DE93",2004,9,"Lüneburg"
"Y20-64","DE94",2004,9.1,"Weser-Ems"
"Y20-64","DEA",2004,9.6,"Nordrhein-Westfalen"
"Y20-64","DEA1",2004,10,"Düsseldorf"
"Y20-64","DEA2",2004,8.4,"Köln"
"Y20-64","DEA3",2004,8.7,"Münster"
"Y20-64","DEA4",2004,9.5,"Detmold"
"Y20-64","DEA5",2004,11,"Arnsberg"
"Y20-64","DEB",2004,7,"Rheinland-Pfalz"
"Y20-64","DEB1",2004,7.6,"Koblenz"
"Y20-64","DEB2",2004,5.9,"Trier"
"Y20-64","DEB3",2004,6.8,"Rheinhessen-Pfalz"
"Y20-64","DEC",2004,8.8,"Saarland"
"Y20-64","DEC0",2004,8.8,"Saarland"
"Y20-64","DED",2004,20,"Sachsen"
"Y20-64","DED2",2004,19.2,"Dresden"
"Y20-64","DEE",2004,23,"Sachsen-Anhalt"
"Y20-64","DEE0",2004,23,"Sachsen-Anhalt"
"Y20-64","DEF",2004,9.7,"Schleswig-Holstein"
"Y20-64","DEF0",2004,9.7,"Schleswig-Holstein"
"Y20-64","DEG",2004,16.9,"Thüringen"
"Y20-64","DEG0",2004,16.9,"Thüringen"
"Y20-64","DK",2004,5.2,"Denmark"
"Y20-64","DK0",2004,5.2,"Danmark"
"Y20-64","EA17",2004,9.1,"Euro area (17 countries)"
"Y20-64","EA18",2004,9.1,"Euro area (18 countries)"
"Y20-64","EA19",2004,9.1,"Euro area (19 countries)"
"Y20-64","EE",2004,9.9,"Estonia"
"Y20-64","EE0",2004,9.9,"Eesti"
"Y20-64","EE00",2004,9.9,"Eesti"
"Y20-64","EL",2004,10.1,"Greece"
"Y20-64","EL1",2004,11.8,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2004,13.1,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2004,11.7,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2004,15.6,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2004,9.7,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2004,10.8,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2004,11,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2004,9.9,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2004,12,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2004,12.3,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2004,8.3,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2004,9.1,"Attiki"
"Y20-64","EL30",2004,9.1,"Attiki"
"Y20-64","EL4",2004,7.2,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2004,9.5,"Voreio Aigaio"
"Y20-64","EL42",2004,8.3,"Notio Aigaio"
"Y20-64","EL43",2004,6,"Kriti"
"Y20-64","ES",2004,10.6,"Spain"
"Y20-64","ES1",2004,12.6,"Noroeste (ES)"
"Y20-64","ES11",2004,14,"Galicia"
"Y20-64","ES12",2004,10,"Principado de Asturias"
"Y20-64","ES13",2004,10.4,"Cantabria"
"Y20-64","ES2",2004,7.4,"Noreste (ES)"
"Y20-64","ES21",2004,9.4,"País Vasco"
"Y20-64","ES22",2004,5.3,"Comunidad Foral de Navarra"
"Y20-64","ES23",2004,5.1,"La Rioja"
"Y20-64","ES24",2004,5.3,"Aragón"
"Y20-64","ES3",2004,6.6,"Comunidad de Madrid"
"Y20-64","ES30",2004,6.6,"Comunidad de Madrid"
"Y20-64","ES4",2004,11.3,"Centro (ES)"
"Y20-64","ES41",2004,10.8,"Castilla y León"
"Y20-64","ES42",2004,8.5,"Castilla-la Mancha"
"Y20-64","ES43",2004,17.7,"Extremadura"
"Y20-64","ES5",2004,9.3,"Este (ES)"
"Y20-64","ES51",2004,9.1,"Cataluña"
"Y20-64","ES52",2004,9.7,"Comunidad Valenciana"
"Y20-64","ES53",2004,8.3,"Illes Balears"
"Y20-64","ES6",2004,15.7,"Sur (ES)"
"Y20-64","ES61",2004,16.8,"Andalucía"
"Y20-64","ES62",2004,10.2,"Región de Murcia"
"Y20-64","ES63",2004,12.2,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2004,17.5,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2004,12.3,"Canarias (ES)"
"Y20-64","ES70",2004,12.3,"Canarias (ES)"
"Y20-64","EU15",2004,8,"European Union (15 countries)"
"Y20-64","EU27",2004,9,"European Union (27 countries)"
"Y20-64","EU28",2004,9,"European Union (28 countries)"
"Y20-64","FI",2004,8.7,"Finland"
"Y20-64","FI1",2004,8.7,"Manner-Suomi"
"Y20-64","FI19",2004,9.3,"Länsi-Suomi"
"Y20-64","FI2",2004,NA,"Åland"
"Y20-64","FI20",2004,NA,"Åland"
"Y20-64","FR",2004,9.1,"France"
"Y20-64","FR1",2004,8.3,"Île de France"
"Y20-64","FR10",2004,8.3,"Île de France"
"Y20-64","FR2",2004,8.4,"Bassin Parisien"
"Y20-64","FR21",2004,8.7,"Champagne-Ardenne"
"Y20-64","FR22",2004,9.8,"Picardie"
"Y20-64","FR23",2004,8.6,"Haute-Normandie"
"Y20-64","FR24",2004,7.1,"Centre (FR)"
"Y20-64","FR25",2004,8.1,"Basse-Normandie"
"Y20-64","FR26",2004,8.4,"Bourgogne"
"Y20-64","FR3",2004,11.8,"Nord - Pas-de-Calais"
"Y20-64","FR30",2004,11.8,"Nord - Pas-de-Calais"
"Y20-64","FR4",2004,9.3,"Est (FR)"
"Y20-64","FR41",2004,11.5,"Lorraine"
"Y20-64","FR42",2004,7.9,"Alsace"
"Y20-64","FR43",2004,7.3,"Franche-Comté"
"Y20-64","FR5",2004,7,"Ouest (FR)"
"Y20-64","FR51",2004,7.6,"Pays de la Loire"
"Y20-64","FR52",2004,6.1,"Bretagne"
"Y20-64","FR53",2004,7.6,"Poitou-Charentes"
"Y20-64","FR6",2004,8.2,"Sud-Ouest (FR)"
"Y20-64","FR61",2004,10.5,"Aquitaine"
"Y20-64","FR62",2004,5.9,"Midi-Pyrénées"
"Y20-64","FR63",2004,NA,"Limousin"
"Y20-64","FR7",2004,8.1,"Centre-Est (FR)"
"Y20-64","FR71",2004,8.1,"Rhône-Alpes"
"Y20-64","FR72",2004,8.1,"Auvergne"
"Y20-64","FR8",2004,10.2,"Méditerranée"
"Y20-64","FR81",2004,10.5,"Languedoc-Roussillon"
"Y20-64","FR82",2004,9.8,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2004,NA,"Corse"
"Y20-64","FR9",2004,26.9,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2004,24.7,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2004,20.9,"Martinique (NUTS 2010)"
"Y20-64","FR93",2004,25.1,"Guyane (NUTS 2010)"
"Y20-64","FR94",2004,31.5,"Réunion (NUTS 2010)"
"Y20-64","HR",2004,13.2,"Croatia"
"Y20-64","HR0",2004,13.2,"Hrvatska"
"Y20-64","HU",2004,5.7,"Hungary"
"Y20-64","HU1",2004,4.1,"Közép-Magyarország"
"Y20-64","HU10",2004,4.1,"Közép-Magyarország"
"Y20-64","HU2",2004,5.3,"Dunántúl"
"Y20-64","HU21",2004,5.2,"Közép-Dunántúl"
"Y20-64","HU22",2004,4.2,"Nyugat-Dunántúl"
"Y20-64","HU23",2004,6.7,"Dél-Dunántúl"
"Y20-64","HU3",2004,7.2,"Alföld és Észak"
"Y20-64","HU31",2004,9.2,"Észak-Magyarország"
"Y20-64","HU32",2004,6.6,"Észak-Alföld"
"Y20-64","HU33",2004,6.1,"Dél-Alföld"
"Y20-64","IE",2004,4.2,"Ireland"
"Y20-64","IE0",2004,4.2,"Éire/Ireland"
"Y20-64","IE01",2004,4.4,"Border, Midland and Western"
"Y20-64","IE02",2004,4.2,"Southern and Eastern"
"Y20-64","IS",2004,3.2,"Iceland"
"Y20-64","IS0",2004,3.2,"Ísland"
"Y20-64","IS00",2004,3.2,"Ísland"
"Y20-64","IT",2004,7.4,"Italy"
"Y20-64","ITC",2004,4,"Nord-Ovest"
"Y20-64","ITC1",2004,5,"Piemonte"
"Y20-64","ITC2",2004,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2004,5.4,"Liguria"
"Y20-64","ITC4",2004,3.4,"Lombardia"
"Y20-64","ITF",2004,13.6,"Sud"
"Y20-64","ITF1",2004,7.3,"Abruzzo"
"Y20-64","ITF2",2004,11.1,"Molise"
"Y20-64","ITF3",2004,14.7,"Campania"
"Y20-64","ITF4",2004,14.9,"Puglia"
"Y20-64","ITF5",2004,11.4,"Basilicata"
"Y20-64","ITF6",2004,13.8,"Calabria"
"Y20-64","ITG",2004,15.5,"Isole"
"Y20-64","ITG1",2004,16.6,"Sicilia"
"Y20-64","ITG2",2004,12.7,"Sardegna"
"Y20-64","ITH",2004,3.5,"Nord-Est"
"Y20-64","ITH1",2004,2.8,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2004,2.4,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2004,3.9,"Veneto"
"Y20-64","ITH4",2004,4,"Friuli-Venezia Giulia"
"Y20-64","ITI",2004,5.8,"Centro (IT)"
"Y20-64","ITI1",2004,5.1,"Toscana"
"Y20-64","ITI2",2004,4.7,"Umbria"
"Y20-64","ITI4",2004,6.8,"Lazio"
"Y20-64","LT",2004,10.5,"Lithuania"
"Y20-64","LT0",2004,10.5,"Lietuva"
"Y20-64","LT00",2004,10.5,"Lietuva"
"Y20-64","LU",2004,4.9,"Luxembourg"
"Y20-64","LU0",2004,4.9,"Luxembourg"
"Y20-64","LU00",2004,4.9,"Luxembourg"
"Y20-64","LV",2004,11.5,"Latvia"
"Y20-64","LV0",2004,11.5,"Latvija"
"Y20-64","LV00",2004,11.5,"Latvija"
"Y20-64","MT",2004,5.5,"Malta"
"Y20-64","MT0",2004,5.5,"Malta"
"Y20-64","MT00",2004,5.5,"Malta"
"Y20-64","NL",2004,4.2,"Netherlands"
"Y20-64","NL1",2004,5.2,"Noord-Nederland"
"Y20-64","NL11",2004,5.6,"Groningen"
"Y20-64","NL12",2004,4.8,"Friesland (NL)"
"Y20-64","NL13",2004,5.2,"Drenthe"
"Y20-64","NL2",2004,4.2,"Oost-Nederland"
"Y20-64","NL21",2004,4.3,"Overijssel"
"Y20-64","NL22",2004,4.1,"Gelderland"
"Y20-64","NL23",2004,4.9,"Flevoland"
"Y20-64","NL3",2004,4,"West-Nederland"
"Y20-64","NL31",2004,3.3,"Utrecht"
"Y20-64","NL32",2004,4.2,"Noord-Holland"
"Y20-64","NL33",2004,4.1,"Zuid-Holland"
"Y20-64","NL34",2004,3.2,"Zeeland"
"Y20-64","NL4",2004,4.2,"Zuid-Nederland"
"Y20-64","NL41",2004,4,"Noord-Brabant"
"Y20-64","NL42",2004,4.5,"Limburg (NL)"
"Y20-64","NO",2004,3.6,"Norway"
"Y20-64","NO0",2004,3.6,"Norge"
"Y20-64","NO01",2004,3.7,"Oslo og Akershus"
"Y20-64","NO02",2004,3.4,"Hedmark og Oppland"
"Y20-64","NO03",2004,3.3,"Sør-Østlandet"
"Y20-64","NO04",2004,4.4,"Agder og Rogaland"
"Y20-64","NO05",2004,3.3,"Vestlandet"
"Y20-64","NO06",2004,3,"Trøndelag"
"Y20-64","NO07",2004,3.7,"Nord-Norge"
"Y20-64","PL",2004,19,"Poland"
"Y20-64","PL1",2004,17,"Region Centralny"
"Y20-64","PL11",2004,18.6,"Lódzkie"
"Y20-64","PL12",2004,16.1,"Mazowieckie"
"Y20-64","PL2",2004,17.7,"Region Poludniowy"
"Y20-64","PL21",2004,16.9,"Malopolskie"
"Y20-64","PL22",2004,18.2,"Slaskie"
"Y20-64","PL3",2004,16.8,"Region Wschodni"
"Y20-64","PL31",2004,16.5,"Lubelskie"
"Y20-64","PL32",2004,15.4,"Podkarpackie"
"Y20-64","PL33",2004,20.9,"Swietokrzyskie"
"Y20-64","PL34",2004,14.9,"Podlaskie"
"Y20-64","PL4",2004,20.1,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2004,17.1,"Wielkopolskie"
"Y20-64","PL42",2004,23.6,"Zachodniopomorskie"
"Y20-64","PL43",2004,24.5,"Lubuskie"
"Y20-64","PL5",2004,24.9,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2004,26.6,"Dolnoslaskie"
"Y20-64","PL52",2004,19,"Opolskie"
"Y20-64","PL6",2004,21.5,"Region Pólnocny"
"Y20-64","PL61",2004,21.9,"Kujawsko-Pomorskie"
"Y20-64","PL62",2004,23.5,"Warminsko-Mazurskie"
"Y20-64","PL63",2004,19.5,"Pomorskie"
"Y20-64","PT",2004,6.4,"Portugal"
"Y20-64","PT1",2004,6.5,"Continente"
"Y20-64","PT11",2004,7.2,"Norte"
"Y20-64","PT15",2004,5.1,"Algarve"
"Y20-64","PT16",2004,4.3,"Centro (PT)"
"Y20-64","PT17",2004,7.3,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2004,8.5,"Alentejo"
"Y20-64","PT2",2004,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2004,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2004,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2004,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2004,7.4,"Romania"
"Y20-64","RO1",2004,6.9,"Macroregiunea unu"
"Y20-64","RO11",2004,5.9,"Nord-Vest"
"Y20-64","RO12",2004,8,"Centru"
"Y20-64","RO2",2004,6.7,"Macroregiunea doi"
"Y20-64","RO21",2004,5.6,"Nord-Est"
"Y20-64","RO22",2004,8.3,"Sud-Est"
"Y20-64","RO3",2004,8.3,"Macroregiunea trei"
"Y20-64","RO31",2004,9.2,"Sud - Muntenia"
"Y20-64","RO32",2004,7.1,"Bucuresti - Ilfov"
"Y20-64","RO4",2004,7.6,"Macroregiunea patru"
"Y20-64","RO41",2004,7.5,"Sud-Vest Oltenia"
"Y20-64","RO42",2004,7.8,"Vest"
"Y20-64","SE",2004,6,"Sweden"
"Y20-64","SE1",2004,5.6,"Östra Sverige"
"Y20-64","SE11",2004,5.2,"Stockholm"
"Y20-64","SE12",2004,6.1,"Östra Mellansverige"
"Y20-64","SE2",2004,6,"Södra Sverige"
"Y20-64","SE21",2004,4.4,"Småland med öarna"
"Y20-64","SE22",2004,7.7,"Sydsverige"
"Y20-64","SE23",2004,5.5,"Västsverige"
"Y20-64","SE3",2004,7,"Norra Sverige"
"Y20-64","SE31",2004,7.5,"Norra Mellansverige"
"Y20-64","SE32",2004,6.2,"Mellersta Norrland"
"Y20-64","SE33",2004,6.6,"Övre Norrland"
"Y20-64","SI",2004,6,"Slovenia"
"Y20-64","SI0",2004,6,"Slovenija"
"Y20-64","SI01",2004,7,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2004,4.8,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2004,18,"Slovakia"
"Y20-64","SK0",2004,18,"Slovensko"
"Y20-64","SK01",2004,8.7,"Bratislavský kraj"
"Y20-64","SK02",2004,13.8,"Západné Slovensko"
"Y20-64","SK03",2004,21.9,"Stredné Slovensko"
"Y20-64","SK04",2004,24.2,"Východné Slovensko"
"Y20-64","UK",2004,4,"United Kingdom"
"Y20-64","UKC",2004,4.5,"North East (UK)"
"Y20-64","UKC1",2004,4.4,"Tees Valley and Durham"
"Y20-64","UKC2",2004,4.7,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2004,3.5,"North West (UK)"
"Y20-64","UKD1",2004,NA,"Cumbria"
"Y20-64","UKD3",2004,3.7,"Greater Manchester"
"Y20-64","UKD4",2004,3.3,"Lancashire"
"Y20-64","UKE",2004,3.6,"Yorkshire and The Humber"
"Y20-64","UKE1",2004,4.2,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2004,NA,"North Yorkshire"
"Y20-64","UKE3",2004,4,"South Yorkshire"
"Y20-64","UKE4",2004,3.7,"West Yorkshire"
"Y20-64","UKF",2004,3.6,"East Midlands (UK)"
"Y20-64","UKF1",2004,3.8,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2004,2.8,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2004,4.7,"Lincolnshire"
"Y20-64","UKG",2004,4.6,"West Midlands (UK)"
"Y20-64","UKG1",2004,2.8,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2004,3.6,"Shropshire and Staffordshire"
"Y20-64","UKG3",2004,6,"West Midlands"
"Y20-64","UKH",2004,3.3,"East of England"
"Y20-64","UKH1",2004,2.9,"East Anglia"
"Y20-64","UKH2",2004,3,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2004,4.1,"Essex"
"Y20-64","UKI",2004,5.8,"London"
"Y20-64","UKI1",2004,8.2,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2004,4.2,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2004,3.2,"South East (UK)"
"Y20-64","UKJ1",2004,3.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2004,2.6,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2004,3.1,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2004,4.2,"Kent"
"Y20-64","UKK",2004,2.5,"South West (UK)"
"Y20-64","UKK1",2004,2.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2004,NA,"Dorset and Somerset"
"Y20-64","UKK3",2004,NA,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2004,3.1,"Devon"
"Y20-64","UKL",2004,3.9,"Wales"
"Y20-64","UKL1",2004,4.5,"West Wales and The Valleys"
"Y20-64","UKL2",2004,3,"East Wales"
"Y20-64","UKM",2004,5.1,"Scotland"
"Y20-64","UKM2",2004,4,"Eastern Scotland"
"Y20-64","UKM3",2004,6.6,"South Western Scotland"
"Y20-64","UKM5",2004,NA,"North Eastern Scotland"
"Y20-64","UKM6",2004,4.3,"Highlands and Islands"
"Y20-64","UKN",2004,4.3,"Northern Ireland (UK)"
"Y20-64","UKN0",2004,4.3,"Northern Ireland (UK)"
"Y_GE15","AT",2004,5.8,"Austria"
"Y_GE15","AT1",2004,7.5,"Ostösterreich"
"Y_GE15","AT11",2004,5.5,"Burgenland (AT)"
"Y_GE15","AT12",2004,4.6,"Niederösterreich"
"Y_GE15","AT13",2004,10.6,"Wien"
"Y_GE15","AT2",2004,5.2,"Südösterreich"
"Y_GE15","AT21",2004,6.3,"Kärnten"
"Y_GE15","AT22",2004,4.7,"Steiermark"
"Y_GE15","AT3",2004,4.3,"Westösterreich"
"Y_GE15","AT31",2004,5,"Oberösterreich"
"Y_GE15","AT32",2004,4.4,"Salzburg"
"Y_GE15","AT33",2004,2.9,"Tirol"
"Y_GE15","AT34",2004,4.2,"Vorarlberg"
"Y_GE15","BE",2004,7.4,"Belgium"
"Y_GE15","BE1",2004,13.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2004,13.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2004,4.5,"Vlaams Gewest"
"Y_GE15","BE21",2004,5.3,"Prov. Antwerpen"
"Y_GE15","BE22",2004,5.9,"Prov. Limburg (BE)"
"Y_GE15","BE23",2004,4.1,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2004,4.4,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2004,3.2,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2004,11,"Région wallonne"
"Y_GE15","BE31",2004,7,"Prov. Brabant Wallon"
"Y_GE15","BE32",2004,12.5,"Prov. Hainaut"
"Y_GE15","BE33",2004,13,"Prov. Liège"
"Y_GE15","BE34",2004,7.1,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2004,7.8,"Prov. Namur"
"Y_GE15","BG",2004,12,"Bulgaria"
"Y_GE15","BG3",2004,14.6,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2004,12.5,"Severozapaden"
"Y_GE15","BG32",2004,14.8,"Severen tsentralen"
"Y_GE15","BG33",2004,17.7,"Severoiztochen"
"Y_GE15","BG34",2004,13.1,"Yugoiztochen"
"Y_GE15","BG4",2004,9.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2004,9.3,"Yugozapaden"
"Y_GE15","BG42",2004,9.7,"Yuzhen tsentralen"
"Y_GE15","CH",2004,4.3,"Switzerland"
"Y_GE15","CH0",2004,4.3,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2004,5.7,"Région lémanique"
"Y_GE15","CH02",2004,3.8,"Espace Mittelland"
"Y_GE15","CH03",2004,3.8,"Nordwestschweiz"
"Y_GE15","CH04",2004,5,"Zürich"
"Y_GE15","CH05",2004,3.5,"Ostschweiz"
"Y_GE15","CH06",2004,3.3,"Zentralschweiz"
"Y_GE15","CH07",2004,5.5,"Ticino"
"Y_GE15","CY",2004,4.3,"Cyprus"
"Y_GE15","CY0",2004,4.3,"Kypros"
"Y_GE15","CY00",2004,4.3,"Kypros"
"Y_GE15","CZ",2004,8.2,"Czech Republic"
"Y_GE15","CZ0",2004,8.2,"Ceská republika"
"Y_GE15","CZ01",2004,3.9,"Praha"
"Y_GE15","CZ02",2004,5.4,"Strední Cechy"
"Y_GE15","CZ03",2004,5.8,"Jihozápad"
"Y_GE15","CZ04",2004,12.1,"Severozápad"
"Y_GE15","CZ05",2004,6.7,"Severovýchod"
"Y_GE15","CZ06",2004,7.9,"Jihovýchod"
"Y_GE15","CZ07",2004,9.9,"Strední Morava"
"Y_GE15","CZ08",2004,14.6,"Moravskoslezsko"
"Y_GE15","DE",2004,10.7,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2004,6.6,"Baden-Württemberg"
"Y_GE15","DE11",2004,6.7,"Stuttgart"
"Y_GE15","DE12",2004,7,"Karlsruhe"
"Y_GE15","DE13",2004,6.4,"Freiburg"
"Y_GE15","DE14",2004,6.2,"Tübingen"
"Y_GE15","DE2",2004,6.8,"Bayern"
"Y_GE15","DE21",2004,5.3,"Oberbayern"
"Y_GE15","DE22",2004,6.4,"Niederbayern"
"Y_GE15","DE23",2004,6.9,"Oberpfalz"
"Y_GE15","DE24",2004,10,"Oberfranken"
"Y_GE15","DE25",2004,8.5,"Mittelfranken"
"Y_GE15","DE26",2004,7.4,"Unterfranken"
"Y_GE15","DE27",2004,6.8,"Schwaben"
"Y_GE15","DE3",2004,19.1,"Berlin"
"Y_GE15","DE30",2004,19.1,"Berlin"
"Y_GE15","DE4",2004,19.2,"Brandenburg"
"Y_GE15","DE40",2004,19.2,"Brandenburg"
"Y_GE15","DE5",2004,14.6,"Bremen"
"Y_GE15","DE50",2004,14.6,"Bremen"
"Y_GE15","DE6",2004,10.6,"Hamburg"
"Y_GE15","DE60",2004,10.6,"Hamburg"
"Y_GE15","DE7",2004,7.9,"Hessen"
"Y_GE15","DE71",2004,7.8,"Darmstadt"
"Y_GE15","DE72",2004,8.5,"Gießen"
"Y_GE15","DE73",2004,7.7,"Kassel"
"Y_GE15","DE8",2004,22.1,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2004,22.1,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2004,9.5,"Niedersachsen"
"Y_GE15","DE91",2004,10.4,"Braunschweig"
"Y_GE15","DE92",2004,9.9,"Hannover"
"Y_GE15","DE93",2004,8.8,"Lüneburg"
"Y_GE15","DE94",2004,9,"Weser-Ems"
"Y_GE15","DEA",2004,9.5,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2004,9.9,"Düsseldorf"
"Y_GE15","DEA2",2004,8.3,"Köln"
"Y_GE15","DEA3",2004,8.7,"Münster"
"Y_GE15","DEA4",2004,9.4,"Detmold"
"Y_GE15","DEA5",2004,10.9,"Arnsberg"
"Y_GE15","DEB",2004,7,"Rheinland-Pfalz"
"Y_GE15","DEB1",2004,7.6,"Koblenz"
"Y_GE15","DEB2",2004,6,"Trier"
"Y_GE15","DEB3",2004,6.9,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2004,8.7,"Saarland"
"Y_GE15","DEC0",2004,8.7,"Saarland"
"Y_GE15","DED",2004,19.4,"Sachsen"
"Y_GE15","DED2",2004,18.7,"Dresden"
"Y_GE15","DEE",2004,22.4,"Sachsen-Anhalt"
"Y_GE15","DEE0",2004,22.4,"Sachsen-Anhalt"
"Y_GE15","DEF",2004,9.7,"Schleswig-Holstein"
"Y_GE15","DEF0",2004,9.7,"Schleswig-Holstein"
"Y_GE15","DEG",2004,16.3,"Thüringen"
"Y_GE15","DEG0",2004,16.3,"Thüringen"
"Y_GE15","DK",2004,5.2,"Denmark"
"Y_GE15","DK0",2004,5.2,"Danmark"
"Y_GE15","EA17",2004,9.3,"Euro area (17 countries)"
"Y_GE15","EA18",2004,9.3,"Euro area (18 countries)"
"Y_GE15","EA19",2004,9.3,"Euro area (19 countries)"
"Y_GE15","EE",2004,10.2,"Estonia"
"Y_GE15","EE0",2004,10.2,"Eesti"
"Y_GE15","EE00",2004,10.2,"Eesti"
"Y_GE15","EL",2004,10.3,"Greece"
"Y_GE15","EL1",2004,12,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2004,13.1,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2004,11.9,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2004,16.3,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2004,9.7,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2004,11.1,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2004,11.5,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2004,10.4,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2004,12.3,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2004,12.4,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2004,8.4,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2004,9.3,"Attiki"
"Y_GE15","EL30",2004,9.3,"Attiki"
"Y_GE15","EL4",2004,7.4,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2004,9.6,"Voreio Aigaio"
"Y_GE15","EL42",2004,8.8,"Notio Aigaio"
"Y_GE15","EL43",2004,6,"Kriti"
"Y_GE15","ES",2004,11.1,"Spain"
"Y_GE15","ES1",2004,12.8,"Noroeste (ES)"
"Y_GE15","ES11",2004,14.1,"Galicia"
"Y_GE15","ES12",2004,10.3,"Principado de Asturias"
"Y_GE15","ES13",2004,10.5,"Cantabria"
"Y_GE15","ES2",2004,7.6,"Noreste (ES)"
"Y_GE15","ES21",2004,9.6,"País Vasco"
"Y_GE15","ES22",2004,5.4,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2004,5.3,"La Rioja"
"Y_GE15","ES24",2004,5.5,"Aragón"
"Y_GE15","ES3",2004,6.9,"Comunidad de Madrid"
"Y_GE15","ES30",2004,6.9,"Comunidad de Madrid"
"Y_GE15","ES4",2004,11.6,"Centro (ES)"
"Y_GE15","ES41",2004,11,"Castilla y León"
"Y_GE15","ES42",2004,8.9,"Castilla-la Mancha"
"Y_GE15","ES43",2004,18,"Extremadura"
"Y_GE15","ES5",2004,9.9,"Este (ES)"
"Y_GE15","ES51",2004,9.8,"Cataluña"
"Y_GE15","ES52",2004,10.3,"Comunidad Valenciana"
"Y_GE15","ES53",2004,9.1,"Illes Balears"
"Y_GE15","ES6",2004,16.3,"Sur (ES)"
"Y_GE15","ES61",2004,17.4,"Andalucía"
"Y_GE15","ES62",2004,10.9,"Región de Murcia"
"Y_GE15","ES63",2004,13.9,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2004,17.3,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2004,12.7,"Canarias (ES)"
"Y_GE15","ES70",2004,12.7,"Canarias (ES)"
"Y_GE15","EU15",2004,8.3,"European Union (15 countries)"
"Y_GE15","EU27",2004,9.2,"European Union (27 countries)"
"Y_GE15","EU28",2004,9.2,"European Union (28 countries)"
"Y_GE15","FI",2004,10.4,"Finland"
"Y_GE15","FI1",2004,10.4,"Manner-Suomi"
"Y_GE15","FI19",2004,11,"Länsi-Suomi"
"Y_GE15","FI2",2004,NA,"Åland"
"Y_GE15","FI20",2004,NA,"Åland"
"Y_GE15","FR",2004,9.4,"France"
"Y_GE15","FR1",2004,8.5,"Île de France"
"Y_GE15","FR10",2004,8.5,"Île de France"
"Y_GE15","FR2",2004,8.8,"Bassin Parisien"
"Y_GE15","FR21",2004,9.2,"Champagne-Ardenne"
"Y_GE15","FR22",2004,10.2,"Picardie"
"Y_GE15","FR23",2004,8.9,"Haute-Normandie"
"Y_GE15","FR24",2004,7.5,"Centre (FR)"
"Y_GE15","FR25",2004,8.7,"Basse-Normandie"
"Y_GE15","FR26",2004,8.6,"Bourgogne"
"Y_GE15","FR3",2004,12.4,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2004,12.4,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2004,9.8,"Est (FR)"
"Y_GE15","FR41",2004,12.3,"Lorraine"
"Y_GE15","FR42",2004,8.3,"Alsace"
"Y_GE15","FR43",2004,7.7,"Franche-Comté"
"Y_GE15","FR5",2004,7.2,"Ouest (FR)"
"Y_GE15","FR51",2004,7.8,"Pays de la Loire"
"Y_GE15","FR52",2004,6.1,"Bretagne"
"Y_GE15","FR53",2004,8,"Poitou-Charentes"
"Y_GE15","FR6",2004,8.4,"Sud-Ouest (FR)"
"Y_GE15","FR61",2004,10.7,"Aquitaine"
"Y_GE15","FR62",2004,6.1,"Midi-Pyrénées"
"Y_GE15","FR63",2004,NA,"Limousin"
"Y_GE15","FR7",2004,8.2,"Centre-Est (FR)"
"Y_GE15","FR71",2004,8.3,"Rhône-Alpes"
"Y_GE15","FR72",2004,8.1,"Auvergne"
"Y_GE15","FR8",2004,10.3,"Méditerranée"
"Y_GE15","FR81",2004,10.9,"Languedoc-Roussillon"
"Y_GE15","FR82",2004,9.9,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2004,NA,"Corse"
"Y_GE15","FR9",2004,27.7,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2004,25.1,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2004,21.5,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2004,25.7,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2004,32.8,"Réunion (NUTS 2010)"
"Y_GE15","HR",2004,13.7,"Croatia"
"Y_GE15","HR0",2004,13.7,"Hrvatska"
"Y_GE15","HU",2004,5.8,"Hungary"
"Y_GE15","HU1",2004,4.2,"Közép-Magyarország"
"Y_GE15","HU10",2004,4.2,"Közép-Magyarország"
"Y_GE15","HU2",2004,5.5,"Dunántúl"
"Y_GE15","HU21",2004,5.3,"Közép-Dunántúl"
"Y_GE15","HU22",2004,4.4,"Nyugat-Dunántúl"
"Y_GE15","HU23",2004,6.9,"Dél-Dunántúl"
"Y_GE15","HU3",2004,7.4,"Alföld és Észak"
"Y_GE15","HU31",2004,9.5,"Észak-Magyarország"
"Y_GE15","HU32",2004,6.8,"Észak-Alföld"
"Y_GE15","HU33",2004,6.2,"Dél-Alföld"
"Y_GE15","IE",2004,4.5,"Ireland"
"Y_GE15","IE0",2004,4.5,"Éire/Ireland"
"Y_GE15","IE01",2004,4.6,"Border, Midland and Western"
"Y_GE15","IE02",2004,4.4,"Southern and Eastern"
"Y_GE15","IS",2004,4,"Iceland"
"Y_GE15","IS0",2004,4,"Ísland"
"Y_GE15","IS00",2004,4,"Ísland"
"Y_GE15","IT",2004,7.9,"Italy"
"Y_GE15","ITC",2004,4.4,"Nord-Ovest"
"Y_GE15","ITC1",2004,5.4,"Piemonte"
"Y_GE15","ITC2",2004,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2004,5.4,"Liguria"
"Y_GE15","ITC4",2004,3.8,"Lombardia"
"Y_GE15","ITF",2004,14.2,"Sud"
"Y_GE15","ITF1",2004,7.9,"Abruzzo"
"Y_GE15","ITF2",2004,11.4,"Molise"
"Y_GE15","ITF3",2004,15.3,"Campania"
"Y_GE15","ITF4",2004,15.3,"Puglia"
"Y_GE15","ITF5",2004,11.6,"Basilicata"
"Y_GE15","ITF6",2004,14.5,"Calabria"
"Y_GE15","ITG",2004,16.1,"Isole"
"Y_GE15","ITG1",2004,17.2,"Sicilia"
"Y_GE15","ITG2",2004,13.4,"Sardegna"
"Y_GE15","ITH",2004,3.9,"Nord-Est"
"Y_GE15","ITH1",2004,3.2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2004,3,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2004,4.3,"Veneto"
"Y_GE15","ITH4",2004,4.3,"Friuli-Venezia Giulia"
"Y_GE15","ITI",2004,6.1,"Centro (IT)"
"Y_GE15","ITI1",2004,5.4,"Toscana"
"Y_GE15","ITI2",2004,5,"Umbria"
"Y_GE15","ITI4",2004,7.2,"Lazio"
"Y_GE15","LT",2004,10.7,"Lithuania"
"Y_GE15","LT0",2004,10.7,"Lietuva"
"Y_GE15","LT00",2004,10.7,"Lietuva"
"Y_GE15","LU",2004,5.1,"Luxembourg"
"Y_GE15","LU0",2004,5.1,"Luxembourg"
"Y_GE15","LU00",2004,5.1,"Luxembourg"
"Y_GE15","LV",2004,11.7,"Latvia"
"Y_GE15","LV0",2004,11.7,"Latvija"
"Y_GE15","LV00",2004,11.7,"Latvija"
"Y_GE15","MT",2004,7.3,"Malta"
"Y_GE15","MT0",2004,7.3,"Malta"
"Y_GE15","MT00",2004,7.3,"Malta"
"Y_GE15","NL",2004,4.6,"Netherlands"
"Y_GE15","NL1",2004,5.6,"Noord-Nederland"
"Y_GE15","NL11",2004,6,"Groningen"
"Y_GE15","NL12",2004,5.2,"Friesland (NL)"
"Y_GE15","NL13",2004,5.5,"Drenthe"
"Y_GE15","NL2",2004,4.7,"Oost-Nederland"
"Y_GE15","NL21",2004,4.7,"Overijssel"
"Y_GE15","NL22",2004,4.4,"Gelderland"
"Y_GE15","NL23",2004,6.5,"Flevoland"
"Y_GE15","NL3",2004,4.4,"West-Nederland"
"Y_GE15","NL31",2004,3.7,"Utrecht"
"Y_GE15","NL32",2004,4.8,"Noord-Holland"
"Y_GE15","NL33",2004,4.5,"Zuid-Holland"
"Y_GE15","NL34",2004,3.3,"Zeeland"
"Y_GE15","NL4",2004,4.6,"Zuid-Nederland"
"Y_GE15","NL41",2004,4.4,"Noord-Brabant"
"Y_GE15","NL42",2004,5,"Limburg (NL)"
"Y_GE15","NO",2004,4.3,"Norway"
"Y_GE15","NO0",2004,4.3,"Norge"
"Y_GE15","NO01",2004,4.2,"Oslo og Akershus"
"Y_GE15","NO02",2004,4.5,"Hedmark og Oppland"
"Y_GE15","NO03",2004,3.9,"Sør-Østlandet"
"Y_GE15","NO04",2004,5,"Agder og Rogaland"
"Y_GE15","NO05",2004,4,"Vestlandet"
"Y_GE15","NO06",2004,3.6,"Trøndelag"
"Y_GE15","NO07",2004,5,"Nord-Norge"
"Y_GE15","PL",2004,19.1,"Poland"
"Y_GE15","PL1",2004,17,"Region Centralny"
"Y_GE15","PL11",2004,18.8,"Lódzkie"
"Y_GE15","PL12",2004,16,"Mazowieckie"
"Y_GE15","PL2",2004,17.8,"Region Poludniowy"
"Y_GE15","PL21",2004,16.8,"Malopolskie"
"Y_GE15","PL22",2004,18.5,"Slaskie"
"Y_GE15","PL3",2004,16.5,"Region Wschodni"
"Y_GE15","PL31",2004,16.1,"Lubelskie"
"Y_GE15","PL32",2004,15.1,"Podkarpackie"
"Y_GE15","PL33",2004,20.4,"Swietokrzyskie"
"Y_GE15","PL34",2004,14.8,"Podlaskie"
"Y_GE15","PL4",2004,20.3,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2004,17.2,"Wielkopolskie"
"Y_GE15","PL42",2004,23.8,"Zachodniopomorskie"
"Y_GE15","PL43",2004,24.9,"Lubuskie"
"Y_GE15","PL5",2004,25,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2004,26.7,"Dolnoslaskie"
"Y_GE15","PL52",2004,19.3,"Opolskie"
"Y_GE15","PL6",2004,21.7,"Region Pólnocny"
"Y_GE15","PL61",2004,22,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2004,23.8,"Warminsko-Mazurskie"
"Y_GE15","PL63",2004,19.8,"Pomorskie"
"Y_GE15","PT",2004,6.3,"Portugal"
"Y_GE15","PT1",2004,6.5,"Continente"
"Y_GE15","PT11",2004,7.3,"Norte"
"Y_GE15","PT15",2004,5,"Algarve"
"Y_GE15","PT16",2004,4,"Centro (PT)"
"Y_GE15","PT17",2004,7.3,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2004,8.8,"Alentejo"
"Y_GE15","PT2",2004,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2004,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2004,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2004,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2004,7.7,"Romania"
"Y_GE15","RO1",2004,7.4,"Macroregiunea unu"
"Y_GE15","RO11",2004,6.2,"Nord-Vest"
"Y_GE15","RO12",2004,8.7,"Centru"
"Y_GE15","RO2",2004,7,"Macroregiunea doi"
"Y_GE15","RO21",2004,5.8,"Nord-Est"
"Y_GE15","RO22",2004,8.7,"Sud-Est"
"Y_GE15","RO3",2004,8.9,"Macroregiunea trei"
"Y_GE15","RO31",2004,9.4,"Sud - Muntenia"
"Y_GE15","RO32",2004,8.2,"Bucuresti - Ilfov"
"Y_GE15","RO4",2004,7.6,"Macroregiunea patru"
"Y_GE15","RO41",2004,7,"Sud-Vest Oltenia"
"Y_GE15","RO42",2004,8.4,"Vest"
"Y_GE15","SE",2004,6.7,"Sweden"
"Y_GE15","SE1",2004,6.2,"Östra Sverige"
"Y_GE15","SE11",2004,5.8,"Stockholm"
"Y_GE15","SE12",2004,6.8,"Östra Mellansverige"
"Y_GE15","SE2",2004,6.7,"Södra Sverige"
"Y_GE15","SE21",2004,5.1,"Småland med öarna"
"Y_GE15","SE22",2004,8.3,"Sydsverige"
"Y_GE15","SE23",2004,6.2,"Västsverige"
"Y_GE15","SE3",2004,7.7,"Norra Sverige"
"Y_GE15","SE31",2004,8.1,"Norra Mellansverige"
"Y_GE15","SE32",2004,7.1,"Mellersta Norrland"
"Y_GE15","SE33",2004,7.5,"Övre Norrland"
"Y_GE15","SI",2004,6,"Slovenia"
"Y_GE15","SI0",2004,6,"Slovenija"
"Y_GE15","SI01",2004,7.1,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2004,4.7,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2004,18.6,"Slovakia"
"Y_GE15","SK0",2004,18.6,"Slovensko"
"Y_GE15","SK01",2004,9.1,"Bratislavský kraj"
"Y_GE15","SK02",2004,14.2,"Západné Slovensko"
"Y_GE15","SK03",2004,22.5,"Stredné Slovensko"
"Y_GE15","SK04",2004,25,"Východné Slovensko"
"Y_GE15","UK",2004,4.6,"United Kingdom"
"Y_GE15","UKC",2004,5.3,"North East (UK)"
"Y_GE15","UKC1",2004,5.3,"Tees Valley and Durham"
"Y_GE15","UKC2",2004,5.3,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2004,4.3,"North West (UK)"
"Y_GE15","UKD1",2004,4.3,"Cumbria"
"Y_GE15","UKD3",2004,4.7,"Greater Manchester"
"Y_GE15","UKD4",2004,4.1,"Lancashire"
"Y_GE15","UKE",2004,4.2,"Yorkshire and The Humber"
"Y_GE15","UKE1",2004,4.5,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2004,2.7,"North Yorkshire"
"Y_GE15","UKE3",2004,4.9,"South Yorkshire"
"Y_GE15","UKE4",2004,4.3,"West Yorkshire"
"Y_GE15","UKF",2004,4,"East Midlands (UK)"
"Y_GE15","UKF1",2004,4,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2004,3.7,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2004,4.7,"Lincolnshire"
"Y_GE15","UKG",2004,5.4,"West Midlands (UK)"
"Y_GE15","UKG1",2004,3.2,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2004,4.3,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2004,7.2,"West Midlands"
"Y_GE15","UKH",2004,3.8,"East of England"
"Y_GE15","UKH1",2004,3.5,"East Anglia"
"Y_GE15","UKH2",2004,3.7,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2004,4.5,"Essex"
"Y_GE15","UKI",2004,6.5,"London"
"Y_GE15","UKI1",2004,9,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2004,4.8,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2004,3.7,"South East (UK)"
"Y_GE15","UKJ1",2004,3.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2004,3,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2004,3.5,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2004,4.7,"Kent"
"Y_GE15","UKK",2004,3.1,"South West (UK)"
"Y_GE15","UKK1",2004,3.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2004,1.8,"Dorset and Somerset"
"Y_GE15","UKK3",2004,4.5,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2004,3.4,"Devon"
"Y_GE15","UKL",2004,4.5,"Wales"
"Y_GE15","UKL1",2004,5.3,"West Wales and The Valleys"
"Y_GE15","UKL2",2004,3.1,"East Wales"
"Y_GE15","UKM",2004,5.9,"Scotland"
"Y_GE15","UKM2",2004,4.7,"Eastern Scotland"
"Y_GE15","UKM3",2004,7.3,"South Western Scotland"
"Y_GE15","UKM5",2004,5.9,"North Eastern Scotland"
"Y_GE15","UKM6",2004,4.7,"Highlands and Islands"
"Y_GE15","UKN",2004,4.7,"Northern Ireland (UK)"
"Y_GE15","UKN0",2004,4.7,"Northern Ireland (UK)"
"Y_GE25","AT",2004,4.8,"Austria"
"Y_GE25","AT1",2004,6.1,"Ostösterreich"
"Y_GE25","AT11",2004,4.3,"Burgenland (AT)"
"Y_GE25","AT12",2004,3.4,"Niederösterreich"
"Y_GE25","AT13",2004,9,"Wien"
"Y_GE25","AT2",2004,4.7,"Südösterreich"
"Y_GE25","AT21",2004,5.6,"Kärnten"
"Y_GE25","AT22",2004,4.3,"Steiermark"
"Y_GE25","AT3",2004,3.3,"Westösterreich"
"Y_GE25","AT31",2004,3.8,"Oberösterreich"
"Y_GE25","AT32",2004,3.4,"Salzburg"
"Y_GE25","AT33",2004,2.3,"Tirol"
"Y_GE25","AT34",2004,3.5,"Vorarlberg"
"Y_GE25","BE",2004,6.3,"Belgium"
"Y_GE25","BE1",2004,13,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2004,13,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2004,3.7,"Vlaams Gewest"
"Y_GE25","BE21",2004,4.2,"Prov. Antwerpen"
"Y_GE25","BE22",2004,4.8,"Prov. Limburg (BE)"
"Y_GE25","BE23",2004,3,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2004,3.6,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2004,3.1,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2004,9.1,"Région wallonne"
"Y_GE25","BE31",2004,5.3,"Prov. Brabant Wallon"
"Y_GE25","BE32",2004,10.2,"Prov. Hainaut"
"Y_GE25","BE33",2004,11.4,"Prov. Liège"
"Y_GE25","BE34",2004,6.1,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2004,6.1,"Prov. Namur"
"Y_GE25","BG",2004,10.8,"Bulgaria"
"Y_GE25","BG3",2004,13.1,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2004,11.6,"Severozapaden"
"Y_GE25","BG32",2004,13.2,"Severen tsentralen"
"Y_GE25","BG33",2004,15.9,"Severoiztochen"
"Y_GE25","BG34",2004,11.5,"Yugoiztochen"
"Y_GE25","BG4",2004,8.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2004,8.4,"Yugozapaden"
"Y_GE25","BG42",2004,8.3,"Yuzhen tsentralen"
"Y_GE25","CH",2004,3.8,"Switzerland"
"Y_GE25","CH0",2004,3.8,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2004,5.1,"Région lémanique"
"Y_GE25","CH02",2004,3.3,"Espace Mittelland"
"Y_GE25","CH03",2004,3.2,"Nordwestschweiz"
"Y_GE25","CH04",2004,4,"Zürich"
"Y_GE25","CH05",2004,3.2,"Ostschweiz"
"Y_GE25","CH06",2004,3.1,"Zentralschweiz"
"Y_GE25","CH07",2004,4.9,"Ticino"
"Y_GE25","CY",2004,3.8,"Cyprus"
"Y_GE25","CY0",2004,3.8,"Kypros"
"Y_GE25","CY00",2004,3.8,"Kypros"
"Y_GE25","CZ",2004,7,"Czech Republic"
"Y_GE25","CZ0",2004,7,"Ceská republika"
"Y_GE25","CZ01",2004,3.6,"Praha"
"Y_GE25","CZ02",2004,5,"Strední Cechy"
"Y_GE25","CZ03",2004,5.2,"Jihozápad"
"Y_GE25","CZ04",2004,10.4,"Severozápad"
"Y_GE25","CZ05",2004,5.7,"Severovýchod"
"Y_GE25","CZ06",2004,6.5,"Jihovýchod"
"Y_GE25","CZ07",2004,8,"Strední Morava"
"Y_GE25","CZ08",2004,12.5,"Moravskoslezsko"
"Y_GE25","DE",2004,10.4,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2004,6.2,"Baden-Württemberg"
"Y_GE25","DE11",2004,6.5,"Stuttgart"
"Y_GE25","DE12",2004,6.7,"Karlsruhe"
"Y_GE25","DE13",2004,5.7,"Freiburg"
"Y_GE25","DE14",2004,5.7,"Tübingen"
"Y_GE25","DE2",2004,6.5,"Bayern"
"Y_GE25","DE21",2004,5,"Oberbayern"
"Y_GE25","DE22",2004,6,"Niederbayern"
"Y_GE25","DE23",2004,7,"Oberpfalz"
"Y_GE25","DE24",2004,9.4,"Oberfranken"
"Y_GE25","DE25",2004,8.6,"Mittelfranken"
"Y_GE25","DE26",2004,6.7,"Unterfranken"
"Y_GE25","DE27",2004,6.5,"Schwaben"
"Y_GE25","DE3",2004,18.8,"Berlin"
"Y_GE25","DE30",2004,18.8,"Berlin"
"Y_GE25","DE4",2004,18.7,"Brandenburg"
"Y_GE25","DE40",2004,18.7,"Brandenburg"
"Y_GE25","DE5",2004,14,"Bremen"
"Y_GE25","DE50",2004,14,"Bremen"
"Y_GE25","DE6",2004,10.2,"Hamburg"
"Y_GE25","DE60",2004,10.2,"Hamburg"
"Y_GE25","DE7",2004,7.4,"Hessen"
"Y_GE25","DE71",2004,7.3,"Darmstadt"
"Y_GE25","DE72",2004,7.9,"Gießen"
"Y_GE25","DE73",2004,7.2,"Kassel"
"Y_GE25","DE8",2004,22.6,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2004,22.6,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2004,9.3,"Niedersachsen"
"Y_GE25","DE91",2004,10.4,"Braunschweig"
"Y_GE25","DE92",2004,9.5,"Hannover"
"Y_GE25","DE93",2004,8.4,"Lüneburg"
"Y_GE25","DE94",2004,8.9,"Weser-Ems"
"Y_GE25","DEA",2004,9.2,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2004,9.7,"Düsseldorf"
"Y_GE25","DEA2",2004,8.2,"Köln"
"Y_GE25","DEA3",2004,8.1,"Münster"
"Y_GE25","DEA4",2004,8.8,"Detmold"
"Y_GE25","DEA5",2004,10.7,"Arnsberg"
"Y_GE25","DEB",2004,6.4,"Rheinland-Pfalz"
"Y_GE25","DEB1",2004,6.8,"Koblenz"
"Y_GE25","DEB2",2004,5.1,"Trier"
"Y_GE25","DEB3",2004,6.3,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2004,8.3,"Saarland"
"Y_GE25","DEC0",2004,8.3,"Saarland"
"Y_GE25","DED",2004,19.7,"Sachsen"
"Y_GE25","DED2",2004,18.9,"Dresden"
"Y_GE25","DEE",2004,23,"Sachsen-Anhalt"
"Y_GE25","DEE0",2004,23,"Sachsen-Anhalt"
"Y_GE25","DEF",2004,9.1,"Schleswig-Holstein"
"Y_GE25","DEF0",2004,9.1,"Schleswig-Holstein"
"Y_GE25","DEG",2004,16.6,"Thüringen"
"Y_GE25","DEG0",2004,16.6,"Thüringen"
"Y_GE25","DK",2004,4.8,"Denmark"
"Y_GE25","DK0",2004,4.8,"Danmark"
"Y_GE25","EA17",2004,8.2,"Euro area (17 countries)"
"Y_GE25","EA18",2004,8.2,"Euro area (18 countries)"
"Y_GE25","EA19",2004,8.2,"Euro area (19 countries)"
"Y_GE25","EE",2004,8.2,"Estonia"
"Y_GE25","EE0",2004,8.2,"Eesti"
"Y_GE25","EE00",2004,8.2,"Eesti"
"Y_GE25","EL",2004,8.5,"Greece"
"Y_GE25","EL1",2004,9.7,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2004,10.9,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2004,9.6,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2004,12.6,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2004,8.1,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2004,9,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2004,8.9,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2004,8.6,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2004,10.4,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2004,10.2,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2004,6.5,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2004,7.8,"Attiki"
"Y_GE25","EL30",2004,7.8,"Attiki"
"Y_GE25","EL4",2004,5.9,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2004,7.9,"Voreio Aigaio"
"Y_GE25","EL42",2004,7.2,"Notio Aigaio"
"Y_GE25","EL43",2004,4.7,"Kriti"
"Y_GE25","ES",2004,9.6,"Spain"
"Y_GE25","ES1",2004,11.1,"Noroeste (ES)"
"Y_GE25","ES11",2004,12.6,"Galicia"
"Y_GE25","ES12",2004,8.2,"Principado de Asturias"
"Y_GE25","ES13",2004,9.3,"Cantabria"
"Y_GE25","ES2",2004,6.4,"Noreste (ES)"
"Y_GE25","ES21",2004,8.1,"País Vasco"
"Y_GE25","ES22",2004,4.7,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2004,4.7,"La Rioja"
"Y_GE25","ES24",2004,4.6,"Aragón"
"Y_GE25","ES3",2004,6.1,"Comunidad de Madrid"
"Y_GE25","ES30",2004,6.1,"Comunidad de Madrid"
"Y_GE25","ES4",2004,10.4,"Centro (ES)"
"Y_GE25","ES41",2004,9.7,"Castilla y León"
"Y_GE25","ES42",2004,7.9,"Castilla-la Mancha"
"Y_GE25","ES43",2004,16.4,"Extremadura"
"Y_GE25","ES5",2004,8.3,"Este (ES)"
"Y_GE25","ES51",2004,8,"Cataluña"
"Y_GE25","ES52",2004,8.9,"Comunidad Valenciana"
"Y_GE25","ES53",2004,7.8,"Illes Balears"
"Y_GE25","ES6",2004,14.4,"Sur (ES)"
"Y_GE25","ES61",2004,15.5,"Andalucía"
"Y_GE25","ES62",2004,9,"Región de Murcia"
"Y_GE25","ES63",2004,8.7,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2004,15.7,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2004,10.6,"Canarias (ES)"
"Y_GE25","ES70",2004,10.6,"Canarias (ES)"
"Y_GE25","EU15",2004,7.2,"European Union (15 countries)"
"Y_GE25","EU27",2004,8,"European Union (27 countries)"
"Y_GE25","EU28",2004,8,"European Union (28 countries)"
"Y_GE25","FI",2004,7.5,"Finland"
"Y_GE25","FI1",2004,7.6,"Manner-Suomi"
"Y_GE25","FI19",2004,8.2,"Länsi-Suomi"
"Y_GE25","FI2",2004,NA,"Åland"
"Y_GE25","FI20",2004,NA,"Åland"
"Y_GE25","FR",2004,8.1,"France"
"Y_GE25","FR1",2004,7.5,"Île de France"
"Y_GE25","FR10",2004,7.5,"Île de France"
"Y_GE25","FR2",2004,7.3,"Bassin Parisien"
"Y_GE25","FR21",2004,7.8,"Champagne-Ardenne"
"Y_GE25","FR22",2004,8.3,"Picardie"
"Y_GE25","FR23",2004,7.7,"Haute-Normandie"
"Y_GE25","FR24",2004,6.3,"Centre (FR)"
"Y_GE25","FR25",2004,7,"Basse-Normandie"
"Y_GE25","FR26",2004,7.5,"Bourgogne"
"Y_GE25","FR3",2004,10,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2004,10,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2004,8.2,"Est (FR)"
"Y_GE25","FR41",2004,10.6,"Lorraine"
"Y_GE25","FR42",2004,6.6,"Alsace"
"Y_GE25","FR43",2004,NA,"Franche-Comté"
"Y_GE25","FR5",2004,6.3,"Ouest (FR)"
"Y_GE25","FR51",2004,7,"Pays de la Loire"
"Y_GE25","FR52",2004,5.5,"Bretagne"
"Y_GE25","FR53",2004,6.1,"Poitou-Charentes"
"Y_GE25","FR6",2004,7.1,"Sud-Ouest (FR)"
"Y_GE25","FR61",2004,9.4,"Aquitaine"
"Y_GE25","FR62",2004,4.9,"Midi-Pyrénées"
"Y_GE25","FR63",2004,NA,"Limousin"
"Y_GE25","FR7",2004,7.4,"Centre-Est (FR)"
"Y_GE25","FR71",2004,7.6,"Rhône-Alpes"
"Y_GE25","FR72",2004,NA,"Auvergne"
"Y_GE25","FR8",2004,9.3,"Méditerranée"
"Y_GE25","FR81",2004,9.6,"Languedoc-Roussillon"
"Y_GE25","FR82",2004,8.9,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2004,NA,"Corse"
"Y_GE25","FR9",2004,24.1,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2004,22.4,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2004,19.2,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2004,23.1,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2004,28.2,"Réunion (NUTS 2010)"
"Y_GE25","HR",2004,11.1,"Croatia"
"Y_GE25","HR0",2004,11.1,"Hrvatska"
"Y_GE25","HU",2004,5,"Hungary"
"Y_GE25","HU1",2004,3.6,"Közép-Magyarország"
"Y_GE25","HU10",2004,3.6,"Közép-Magyarország"
"Y_GE25","HU2",2004,4.8,"Dunántúl"
"Y_GE25","HU21",2004,4.7,"Közép-Dunántúl"
"Y_GE25","HU22",2004,3.9,"Nyugat-Dunántúl"
"Y_GE25","HU23",2004,5.9,"Dél-Dunántúl"
"Y_GE25","HU3",2004,6.4,"Alföld és Észak"
"Y_GE25","HU31",2004,8.4,"Észak-Magyarország"
"Y_GE25","HU32",2004,5.9,"Észak-Alföld"
"Y_GE25","HU33",2004,5.3,"Dél-Alföld"
"Y_GE25","IE",2004,3.8,"Ireland"
"Y_GE25","IE0",2004,3.8,"Éire/Ireland"
"Y_GE25","IE01",2004,3.9,"Border, Midland and Western"
"Y_GE25","IE02",2004,3.7,"Southern and Eastern"
"Y_GE25","IS",2004,2.3,"Iceland"
"Y_GE25","IS0",2004,2.3,"Ísland"
"Y_GE25","IS00",2004,2.3,"Ísland"
"Y_GE25","IT",2004,6.2,"Italy"
"Y_GE25","ITC",2004,3.6,"Nord-Ovest"
"Y_GE25","ITC1",2004,4.5,"Piemonte"
"Y_GE25","ITC2",2004,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2004,4.6,"Liguria"
"Y_GE25","ITC4",2004,3,"Lombardia"
"Y_GE25","ITF",2004,11.3,"Sud"
"Y_GE25","ITF1",2004,6,"Abruzzo"
"Y_GE25","ITF2",2004,9.3,"Molise"
"Y_GE25","ITF3",2004,12.1,"Campania"
"Y_GE25","ITF4",2004,12.7,"Puglia"
"Y_GE25","ITF5",2004,9.6,"Basilicata"
"Y_GE25","ITF6",2004,11,"Calabria"
"Y_GE25","ITG",2004,13,"Isole"
"Y_GE25","ITG1",2004,14,"Sicilia"
"Y_GE25","ITG2",2004,10.3,"Sardegna"
"Y_GE25","ITH",2004,3,"Nord-Est"
"Y_GE25","ITH1",2004,2.7,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2004,1.9,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2004,3.5,"Veneto"
"Y_GE25","ITH4",2004,3.5,"Friuli-Venezia Giulia"
"Y_GE25","ITI",2004,4.7,"Centro (IT)"
"Y_GE25","ITI1",2004,4.4,"Toscana"
"Y_GE25","ITI2",2004,4.1,"Umbria"
"Y_GE25","ITI4",2004,5.4,"Lazio"
"Y_GE25","LT",2004,9.8,"Lithuania"
"Y_GE25","LT0",2004,9.8,"Lietuva"
"Y_GE25","LT00",2004,9.8,"Lietuva"
"Y_GE25","LU",2004,4.2,"Luxembourg"
"Y_GE25","LU0",2004,4.2,"Luxembourg"
"Y_GE25","LU00",2004,4.2,"Luxembourg"
"Y_GE25","LV",2004,10.4,"Latvia"
"Y_GE25","LV0",2004,10.4,"Latvija"
"Y_GE25","LV00",2004,10.4,"Latvija"
"Y_GE25","MT",2004,4.4,"Malta"
"Y_GE25","MT0",2004,4.4,"Malta"
"Y_GE25","MT00",2004,4.4,"Malta"
"Y_GE25","NL",2004,4,"Netherlands"
"Y_GE25","NL1",2004,4.9,"Noord-Nederland"
"Y_GE25","NL11",2004,5.4,"Groningen"
"Y_GE25","NL12",2004,4.7,"Friesland (NL)"
"Y_GE25","NL13",2004,4.6,"Drenthe"
"Y_GE25","NL2",2004,3.9,"Oost-Nederland"
"Y_GE25","NL21",2004,3.7,"Overijssel"
"Y_GE25","NL22",2004,3.9,"Gelderland"
"Y_GE25","NL23",2004,4.5,"Flevoland"
"Y_GE25","NL3",2004,3.8,"West-Nederland"
"Y_GE25","NL31",2004,3,"Utrecht"
"Y_GE25","NL32",2004,3.9,"Noord-Holland"
"Y_GE25","NL33",2004,4,"Zuid-Holland"
"Y_GE25","NL34",2004,3,"Zeeland"
"Y_GE25","NL4",2004,4.1,"Zuid-Nederland"
"Y_GE25","NL41",2004,3.9,"Noord-Brabant"
"Y_GE25","NL42",2004,4.5,"Limburg (NL)"
"Y_GE25","NO",2004,2.9,"Norway"
"Y_GE25","NO0",2004,2.9,"Norge"
"Y_GE25","NO01",2004,3.1,"Oslo og Akershus"
"Y_GE25","NO02",2004,2.9,"Hedmark og Oppland"
"Y_GE25","NO03",2004,2.4,"Sør-Østlandet"
"Y_GE25","NO04",2004,3.6,"Agder og Rogaland"
"Y_GE25","NO05",2004,2.7,"Vestlandet"
"Y_GE25","NO06",2004,2.5,"Trøndelag"
"Y_GE25","NO07",2004,2.8,"Nord-Norge"
"Y_GE25","PL",2004,16.1,"Poland"
"Y_GE25","PL1",2004,14.5,"Region Centralny"
"Y_GE25","PL11",2004,16.2,"Lódzkie"
"Y_GE25","PL12",2004,13.6,"Mazowieckie"
"Y_GE25","PL2",2004,14.3,"Region Poludniowy"
"Y_GE25","PL21",2004,13.6,"Malopolskie"
"Y_GE25","PL22",2004,14.8,"Slaskie"
"Y_GE25","PL3",2004,13.8,"Region Wschodni"
"Y_GE25","PL31",2004,13.5,"Lubelskie"
"Y_GE25","PL32",2004,12.5,"Podkarpackie"
"Y_GE25","PL33",2004,17.8,"Swietokrzyskie"
"Y_GE25","PL34",2004,12.2,"Podlaskie"
"Y_GE25","PL4",2004,17,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2004,13.9,"Wielkopolskie"
"Y_GE25","PL42",2004,21.4,"Zachodniopomorskie"
"Y_GE25","PL43",2004,20.5,"Lubuskie"
"Y_GE25","PL5",2004,21.6,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2004,23.2,"Dolnoslaskie"
"Y_GE25","PL52",2004,16.3,"Opolskie"
"Y_GE25","PL6",2004,19,"Region Pólnocny"
"Y_GE25","PL61",2004,19.1,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2004,20.8,"Warminsko-Mazurskie"
"Y_GE25","PL63",2004,17.5,"Pomorskie"
"Y_GE25","PT",2004,5.4,"Portugal"
"Y_GE25","PT1",2004,5.6,"Continente"
"Y_GE25","PT11",2004,6.3,"Norte"
"Y_GE25","PT15",2004,4.3,"Algarve"
"Y_GE25","PT16",2004,3.5,"Centro (PT)"
"Y_GE25","PT17",2004,6.3,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2004,7,"Alentejo"
"Y_GE25","PT2",2004,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2004,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2004,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2004,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2004,5.7,"Romania"
"Y_GE25","RO1",2004,5.4,"Macroregiunea unu"
"Y_GE25","RO11",2004,4.4,"Nord-Vest"
"Y_GE25","RO12",2004,6.4,"Centru"
"Y_GE25","RO2",2004,5.3,"Macroregiunea doi"
"Y_GE25","RO21",2004,4.1,"Nord-Est"
"Y_GE25","RO22",2004,6.9,"Sud-Est"
"Y_GE25","RO3",2004,6.5,"Macroregiunea trei"
"Y_GE25","RO31",2004,6.8,"Sud - Muntenia"
"Y_GE25","RO32",2004,6,"Bucuresti - Ilfov"
"Y_GE25","RO4",2004,6,"Macroregiunea patru"
"Y_GE25","RO41",2004,5.9,"Sud-Vest Oltenia"
"Y_GE25","RO42",2004,6,"Vest"
"Y_GE25","SE",2004,5.2,"Sweden"
"Y_GE25","SE1",2004,4.7,"Östra Sverige"
"Y_GE25","SE11",2004,4.4,"Stockholm"
"Y_GE25","SE12",2004,5.1,"Östra Mellansverige"
"Y_GE25","SE2",2004,5.2,"Södra Sverige"
"Y_GE25","SE21",2004,3.7,"Småland med öarna"
"Y_GE25","SE22",2004,6.7,"Sydsverige"
"Y_GE25","SE23",2004,4.8,"Västsverige"
"Y_GE25","SE3",2004,6.1,"Norra Sverige"
"Y_GE25","SE31",2004,6.6,"Norra Mellansverige"
"Y_GE25","SE32",2004,5.3,"Mellersta Norrland"
"Y_GE25","SE33",2004,6,"Övre Norrland"
"Y_GE25","SI",2004,5,"Slovenia"
"Y_GE25","SI0",2004,5,"Slovenija"
"Y_GE25","SI01",2004,5.9,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2004,4.1,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2004,16.4,"Slovakia"
"Y_GE25","SK0",2004,16.4,"Slovensko"
"Y_GE25","SK01",2004,7.6,"Bratislavský kraj"
"Y_GE25","SK02",2004,12.7,"Západné Slovensko"
"Y_GE25","SK03",2004,20.2,"Stredné Slovensko"
"Y_GE25","SK04",2004,22,"Východné Slovensko"
"Y_GE25","UK",2004,3.5,"United Kingdom"
"Y_GE25","UKC",2004,3.8,"North East (UK)"
"Y_GE25","UKC1",2004,3.7,"Tees Valley and Durham"
"Y_GE25","UKC2",2004,3.9,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2004,3,"North West (UK)"
"Y_GE25","UKD1",2004,NA,"Cumbria"
"Y_GE25","UKD3",2004,3,"Greater Manchester"
"Y_GE25","UKD4",2004,3,"Lancashire"
"Y_GE25","UKE",2004,3.3,"Yorkshire and The Humber"
"Y_GE25","UKE1",2004,3.9,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2004,NA,"North Yorkshire"
"Y_GE25","UKE3",2004,3.9,"South Yorkshire"
"Y_GE25","UKE4",2004,3.3,"West Yorkshire"
"Y_GE25","UKF",2004,3.3,"East Midlands (UK)"
"Y_GE25","UKF1",2004,3.5,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2004,2.7,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2004,4.2,"Lincolnshire"
"Y_GE25","UKG",2004,4,"West Midlands (UK)"
"Y_GE25","UKG1",2004,2.5,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2004,3.5,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2004,5.3,"West Midlands"
"Y_GE25","UKH",2004,2.8,"East of England"
"Y_GE25","UKH1",2004,2.3,"East Anglia"
"Y_GE25","UKH2",2004,2.8,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2004,3.6,"Essex"
"Y_GE25","UKI",2004,5.1,"London"
"Y_GE25","UKI1",2004,7.2,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2004,3.7,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2004,2.9,"South East (UK)"
"Y_GE25","UKJ1",2004,3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2004,2.3,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2004,2.7,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2004,3.9,"Kent"
"Y_GE25","UKK",2004,2.4,"South West (UK)"
"Y_GE25","UKK1",2004,2.6,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2004,NA,"Dorset and Somerset"
"Y_GE25","UKK3",2004,NA,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2004,2.7,"Devon"
"Y_GE25","UKL",2004,3.2,"Wales"
"Y_GE25","UKL1",2004,3.8,"West Wales and The Valleys"
"Y_GE25","UKL2",2004,2.3,"East Wales"
"Y_GE25","UKM",2004,4.5,"Scotland"
"Y_GE25","UKM2",2004,3.3,"Eastern Scotland"
"Y_GE25","UKM3",2004,5.9,"South Western Scotland"
"Y_GE25","UKM5",2004,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2004,4.4,"Highlands and Islands"
"Y_GE25","UKN",2004,3.7,"Northern Ireland (UK)"
"Y_GE25","UKN0",2004,3.7,"Northern Ireland (UK)"
"Y15-24","AT",2003,7.5,"Austria"
"Y15-24","AT1",2003,10.1,"Ostösterreich"
"Y15-24","AT11",2003,NA,"Burgenland (AT)"
"Y15-24","AT12",2003,6,"Niederösterreich"
"Y15-24","AT13",2003,15,"Wien"
"Y15-24","AT2",2003,6.4,"Südösterreich"
"Y15-24","AT21",2003,NA,"Kärnten"
"Y15-24","AT22",2003,5.5,"Steiermark"
"Y15-24","AT3",2003,5.6,"Westösterreich"
"Y15-24","AT31",2003,6.4,"Oberösterreich"
"Y15-24","AT32",2003,NA,"Salzburg"
"Y15-24","AT33",2003,NA,"Tirol"
"Y15-24","AT34",2003,NA,"Vorarlberg"
"Y15-24","BE",2003,19,"Belgium"
"Y15-24","BE1",2003,35.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2003,35.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2003,13.5,"Vlaams Gewest"
"Y15-24","BE21",2003,15.9,"Prov. Antwerpen"
"Y15-24","BE22",2003,14.5,"Prov. Limburg (BE)"
"Y15-24","BE23",2003,13.6,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2003,15.2,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2003,9.1,"Prov. West-Vlaanderen"
"Y15-24","BE3",2003,26.2,"Région wallonne"
"Y15-24","BE31",2003,NA,"Prov. Brabant Wallon"
"Y15-24","BE32",2003,35.6,"Prov. Hainaut"
"Y15-24","BE33",2003,20.6,"Prov. Liège"
"Y15-24","BE34",2003,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2003,NA,"Prov. Namur"
"Y15-24","BG",2003,27.1,"Bulgaria"
"Y15-24","BG3",2003,30.8,"Severna i yugoiztochna Bulgaria"
"Y15-24","BG31",2003,27,"Severozapaden"
"Y15-24","BG32",2003,29.5,"Severen tsentralen"
"Y15-24","BG33",2003,30.7,"Severoiztochen"
"Y15-24","BG34",2003,34.4,"Yugoiztochen"
"Y15-24","BG4",2003,23.1,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y15-24","BG41",2003,21,"Yugozapaden"
"Y15-24","BG42",2003,26.2,"Yuzhen tsentralen"
"Y15-24","CH",2003,8.5,"Switzerland"
"Y15-24","CH0",2003,8.5,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2003,11.9,"Région lémanique"
"Y15-24","CH02",2003,8.5,"Espace Mittelland"
"Y15-24","CH03",2003,7,"Nordwestschweiz"
"Y15-24","CH04",2003,7.1,"Zürich"
"Y15-24","CH05",2003,7.5,"Ostschweiz"
"Y15-24","CH06",2003,7.8,"Zentralschweiz"
"Y15-24","CH07",2003,12.1,"Ticino"
"Y15-24","CY",2003,8.9,"Cyprus"
"Y15-24","CY0",2003,8.9,"Kypros"
"Y15-24","CY00",2003,8.9,"Kypros"
"Y15-24","CZ",2003,16.8,"Czech Republic"
"Y15-24","CZ0",2003,16.8,"Ceská republika"
"Y15-24","CZ01",2003,10.5,"Praha"
"Y15-24","CZ02",2003,6,"Strední Cechy"
"Y15-24","CZ03",2003,11.6,"Jihozápad"
"Y15-24","CZ04",2003,19.7,"Severozápad"
"Y15-24","CZ05",2003,16.2,"Severovýchod"
"Y15-24","CZ06",2003,18.2,"Jihovýchod"
"Y15-24","CZ07",2003,19.9,"Strední Morava"
"Y15-24","CZ08",2003,28.8,"Moravskoslezsko"
"Y15-24","DE",2003,11,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2003,7.4,"Baden-Württemberg"
"Y15-24","DE11",2003,8.2,"Stuttgart"
"Y15-24","DE12",2003,7,"Karlsruhe"
"Y15-24","DE13",2003,6,"Freiburg"
"Y15-24","DE14",2003,8,"Tübingen"
"Y15-24","DE2",2003,7.2,"Bayern"
"Y15-24","DE21",2003,6.3,"Oberbayern"
"Y15-24","DE22",2003,7.5,"Niederbayern"
"Y15-24","DE23",2003,7,"Oberpfalz"
"Y15-24","DE24",2003,10.7,"Oberfranken"
"Y15-24","DE25",2003,5.8,"Mittelfranken"
"Y15-24","DE26",2003,8.2,"Unterfranken"
"Y15-24","DE27",2003,7.3,"Schwaben"
"Y15-24","DE3",2003,21.4,"Berlin"
"Y15-24","DE30",2003,21.4,"Berlin"
"Y15-24","DE4",2003,19.4,"Brandenburg"
"Y15-24","DE40",2003,19.4,"Brandenburg"
"Y15-24","DE5",2003,16.6,"Bremen"
"Y15-24","DE50",2003,16.6,"Bremen"
"Y15-24","DE6",2003,9.2,"Hamburg"
"Y15-24","DE60",2003,9.2,"Hamburg"
"Y15-24","DE7",2003,10.6,"Hessen"
"Y15-24","DE71",2003,9.8,"Darmstadt"
"Y15-24","DE72",2003,11.1,"Gießen"
"Y15-24","DE73",2003,12.3,"Kassel"
"Y15-24","DE8",2003,19.8,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2003,19.8,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2003,9.9,"Niedersachsen"
"Y15-24","DE91",2003,13.3,"Braunschweig"
"Y15-24","DE92",2003,7.9,"Hannover"
"Y15-24","DE93",2003,10.3,"Lüneburg"
"Y15-24","DE94",2003,9.2,"Weser-Ems"
"Y15-24","DEA",2003,10.7,"Nordrhein-Westfalen"
"Y15-24","DEA1",2003,12.5,"Düsseldorf"
"Y15-24","DEA2",2003,12.1,"Köln"
"Y15-24","DEA3",2003,9.7,"Münster"
"Y15-24","DEA4",2003,10.3,"Detmold"
"Y15-24","DEA5",2003,7.9,"Arnsberg"
"Y15-24","DEB",2003,7,"Rheinland-Pfalz"
"Y15-24","DEB1",2003,9.8,"Koblenz"
"Y15-24","DEB2",2003,NA,"Trier"
"Y15-24","DEB3",2003,5.8,"Rheinhessen-Pfalz"
"Y15-24","DEC",2003,10.9,"Saarland"
"Y15-24","DEC0",2003,10.9,"Saarland"
"Y15-24","DED",2003,16.6,"Sachsen"
"Y15-24","DED2",2003,17.6,"Dresden"
"Y15-24","DEE",2003,15.2,"Sachsen-Anhalt"
"Y15-24","DEE0",2003,15.2,"Sachsen-Anhalt"
"Y15-24","DEF",2003,9.7,"Schleswig-Holstein"
"Y15-24","DEF0",2003,9.7,"Schleswig-Holstein"
"Y15-24","DEG",2003,12.4,"Thüringen"
"Y15-24","DEG0",2003,12.4,"Thüringen"
"Y15-24","DK",2003,9.8,"Denmark"
"Y15-24","DK0",2003,9.8,"Danmark"
"Y15-24","EA17",2003,17.1,"Euro area (17 countries)"
"Y15-24","EA18",2003,17.1,"Euro area (18 countries)"
"Y15-24","EA19",2003,17.2,"Euro area (19 countries)"
"Y15-24","EE",2003,26.9,"Estonia"
"Y15-24","EE0",2003,26.9,"Eesti"
"Y15-24","EE00",2003,26.9,"Eesti"
"Y15-24","EL",2003,25.4,"Greece"
"Y15-24","EL1",2003,26.7,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2003,22.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2003,25.1,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2003,41.2,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2003,28.6,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2003,28.4,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2003,34.6,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2003,31.5,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2003,30.2,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2003,22,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2003,28,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2003,23.8,"Attiki"
"Y15-24","EL30",2003,23.8,"Attiki"
"Y15-24","EL4",2003,22.2,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2003,31.7,"Voreio Aigaio"
"Y15-24","EL42",2003,21.8,"Notio Aigaio"
"Y15-24","EL43",2003,20.1,"Kriti"
"Y15-24","ES",2003,22.3,"Spain"
"Y15-24","ES1",2003,23.6,"Noroeste (ES)"
"Y15-24","ES11",2003,24.4,"Galicia"
"Y15-24","ES12",2003,24.2,"Principado de Asturias"
"Y15-24","ES13",2003,18.8,"Cantabria"
"Y15-24","ES2",2003,18.5,"Noreste (ES)"
"Y15-24","ES21",2003,23.2,"País Vasco"
"Y15-24","ES22",2003,14.3,"Comunidad Foral de Navarra"
"Y15-24","ES23",2003,NA,"La Rioja"
"Y15-24","ES24",2003,15.1,"Aragón"
"Y15-24","ES3",2003,14.3,"Comunidad de Madrid"
"Y15-24","ES30",2003,14.3,"Comunidad de Madrid"
"Y15-24","ES4",2003,20.8,"Centro (ES)"
"Y15-24","ES41",2003,24.9,"Castilla y León"
"Y15-24","ES42",2003,16.4,"Castilla-la Mancha"
"Y15-24","ES43",2003,21.4,"Extremadura"
"Y15-24","ES5",2003,22.5,"Este (ES)"
"Y15-24","ES51",2003,23.9,"Cataluña"
"Y15-24","ES52",2003,20.2,"Comunidad Valenciana"
"Y15-24","ES53",2003,24.2,"Illes Balears"
"Y15-24","ES6",2003,27.3,"Sur (ES)"
"Y15-24","ES61",2003,29.5,"Andalucía"
"Y15-24","ES62",2003,17.1,"Región de Murcia"
"Y15-24","ES63",2003,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2003,NA,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2003,24,"Canarias (ES)"
"Y15-24","ES70",2003,24,"Canarias (ES)"
"Y15-24","EU15",2003,15.5,"European Union (15 countries)"
"Y15-24","EU27",2003,18.2,"European Union (27 countries)"
"Y15-24","EU28",2003,18.3,"European Union (28 countries)"
"Y15-24","FI",2003,27.8,"Finland"
"Y15-24","FI1",2003,27.9,"Manner-Suomi"
"Y15-24","FI19",2003,28,"Länsi-Suomi"
"Y15-24","FI2",2003,NA,"Åland"
"Y15-24","FI20",2003,NA,"Åland"
"Y15-24","FR",2003,18.2,"France"
"Y15-24","FR1",2003,16.7,"Île de France"
"Y15-24","FR10",2003,16.7,"Île de France"
"Y15-24","FR2",2003,15.2,"Bassin Parisien"
"Y15-24","FR21",2003,NA,"Champagne-Ardenne"
"Y15-24","FR22",2003,NA,"Picardie"
"Y15-24","FR23",2003,NA,"Haute-Normandie"
"Y15-24","FR24",2003,NA,"Centre (FR)"
"Y15-24","FR25",2003,NA,"Basse-Normandie"
"Y15-24","FR26",2003,NA,"Bourgogne"
"Y15-24","FR3",2003,20.8,"Nord - Pas-de-Calais"
"Y15-24","FR30",2003,20.8,"Nord - Pas-de-Calais"
"Y15-24","FR4",2003,22.3,"Est (FR)"
"Y15-24","FR41",2003,NA,"Lorraine"
"Y15-24","FR42",2003,NA,"Alsace"
"Y15-24","FR43",2003,NA,"Franche-Comté"
"Y15-24","FR5",2003,14.5,"Ouest (FR)"
"Y15-24","FR51",2003,NA,"Pays de la Loire"
"Y15-24","FR52",2003,NA,"Bretagne"
"Y15-24","FR53",2003,NA,"Poitou-Charentes"
"Y15-24","FR6",2003,19.6,"Sud-Ouest (FR)"
"Y15-24","FR61",2003,NA,"Aquitaine"
"Y15-24","FR62",2003,NA,"Midi-Pyrénées"
"Y15-24","FR63",2003,NA,"Limousin"
"Y15-24","FR7",2003,12,"Centre-Est (FR)"
"Y15-24","FR71",2003,12.5,"Rhône-Alpes"
"Y15-24","FR72",2003,NA,"Auvergne"
"Y15-24","FR8",2003,22.3,"Méditerranée"
"Y15-24","FR81",2003,NA,"Languedoc-Roussillon"
"Y15-24","FR82",2003,19.4,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2003,NA,"Corse"
"Y15-24","FR9",2003,52.6,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2003,56,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2003,48.7,"Martinique (NUTS 2010)"
"Y15-24","FR93",2003,49.8,"Guyane (NUTS 2010)"
"Y15-24","FR94",2003,53,"Réunion (NUTS 2010)"
"Y15-24","HR",2003,35.8,"Croatia"
"Y15-24","HR0",2003,35.8,"Hrvatska"
"Y15-24","HU",2003,12.9,"Hungary"
"Y15-24","HU1",2003,10.1,"Közép-Magyarország"
"Y15-24","HU10",2003,10.1,"Közép-Magyarország"
"Y15-24","HU2",2003,12.1,"Dunántúl"
"Y15-24","HU21",2003,9.9,"Közép-Dunántúl"
"Y15-24","HU22",2003,11,"Nyugat-Dunántúl"
"Y15-24","HU23",2003,16.2,"Dél-Dunántúl"
"Y15-24","HU3",2003,15.5,"Alföld és Észak"
"Y15-24","HU31",2003,20.6,"Észak-Magyarország"
"Y15-24","HU32",2003,13,"Észak-Alföld"
"Y15-24","HU33",2003,13.3,"Dél-Alföld"
"Y15-24","IE",2003,8.1,"Ireland"
"Y15-24","IE0",2003,8.1,"Éire/Ireland"
"Y15-24","IE01",2003,10.4,"Border, Midland and Western"
"Y15-24","IE02",2003,7.4,"Southern and Eastern"
"Y15-24","IS",2003,12.5,"Iceland"
"Y15-24","IS0",2003,12.5,"Ísland"
"Y15-24","IS00",2003,12.5,"Ísland"
"Y15-24","IT",2003,26.8,"Italy"
"Y15-24","ITC",2003,12.4,"Nord-Ovest"
"Y15-24","ITC1",2003,16.5,"Piemonte"
"Y15-24","ITC2",2003,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2003,21.3,"Liguria"
"Y15-24","ITC4",2003,9.8,"Lombardia"
"Y15-24","ITF",2003,48.8,"Sud"
"Y15-24","ITF1",2003,12.8,"Abruzzo"
"Y15-24","ITF2",2003,43,"Molise"
"Y15-24","ITF3",2003,59.6,"Campania"
"Y15-24","ITF4",2003,38.9,"Puglia"
"Y15-24","ITF5",2003,41.8,"Basilicata"
"Y15-24","ITF6",2003,55.1,"Calabria"
"Y15-24","ITG",2003,50.4,"Isole"
"Y15-24","ITG1",2003,52.8,"Sicilia"
"Y15-24","ITG2",2003,43.5,"Sardegna"
"Y15-24","ITH",2003,7.2,"Nord-Est"
"Y15-24","ITH1",2003,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2003,NA,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2003,6.8,"Veneto"
"Y15-24","ITH4",2003,14.3,"Friuli-Venezia Giulia"
"Y15-24","ITI",2003,23.4,"Centro (IT)"
"Y15-24","ITI1",2003,14.4,"Toscana"
"Y15-24","ITI2",2003,17.5,"Umbria"
"Y15-24","ITI4",2003,35.1,"Lazio"
"Y15-24","LT",2003,26.9,"Lithuania"
"Y15-24","LT0",2003,26.9,"Lietuva"
"Y15-24","LT00",2003,26.9,"Lietuva"
"Y15-24","LU",2003,10.9,"Luxembourg"
"Y15-24","LU0",2003,10.9,"Luxembourg"
"Y15-24","LU00",2003,10.9,"Luxembourg"
"Y15-24","LV",2003,20.4,"Latvia"
"Y15-24","LV0",2003,20.4,"Latvija"
"Y15-24","LV00",2003,20.4,"Latvija"
"Y15-24","MT",2003,17.4,"Malta"
"Y15-24","MT0",2003,17.4,"Malta"
"Y15-24","MT00",2003,17.4,"Malta"
"Y15-24","NL",2003,6.6,"Netherlands"
"Y15-24","NL1",2003,6.6,"Noord-Nederland"
"Y15-24","NL11",2003,6.9,"Groningen"
"Y15-24","NL12",2003,5.9,"Friesland (NL)"
"Y15-24","NL13",2003,7,"Drenthe"
"Y15-24","NL2",2003,6.1,"Oost-Nederland"
"Y15-24","NL21",2003,5.7,"Overijssel"
"Y15-24","NL22",2003,6.3,"Gelderland"
"Y15-24","NL23",2003,6.1,"Flevoland"
"Y15-24","NL3",2003,7.1,"West-Nederland"
"Y15-24","NL31",2003,6.9,"Utrecht"
"Y15-24","NL32",2003,8.2,"Noord-Holland"
"Y15-24","NL33",2003,6.8,"Zuid-Holland"
"Y15-24","NL34",2003,NA,"Zeeland"
"Y15-24","NL4",2003,6.1,"Zuid-Nederland"
"Y15-24","NL41",2003,6.2,"Noord-Brabant"
"Y15-24","NL42",2003,5.9,"Limburg (NL)"
"Y15-24","NO",2003,11.9,"Norway"
"Y15-24","NO0",2003,11.9,"Norge"
"Y15-24","NO01",2003,9,"Oslo og Akershus"
"Y15-24","NO02",2003,10.7,"Hedmark og Oppland"
"Y15-24","NO03",2003,14.2,"Sør-Østlandet"
"Y15-24","NO04",2003,8.9,"Agder og Rogaland"
"Y15-24","NO05",2003,13.2,"Vestlandet"
"Y15-24","NO06",2003,10.3,"Trøndelag"
"Y15-24","NO07",2003,16.6,"Nord-Norge"
"Y15-24","PL",2003,41.4,"Poland"
"Y15-24","PL1",2003,37.4,"Region Centralny"
"Y15-24","PL11",2003,39.2,"Lódzkie"
"Y15-24","PL12",2003,36.3,"Mazowieckie"
"Y15-24","PL2",2003,44.7,"Region Poludniowy"
"Y15-24","PL21",2003,40,"Malopolskie"
"Y15-24","PL22",2003,49.1,"Slaskie"
"Y15-24","PL3",2003,38.1,"Region Wschodni"
"Y15-24","PL31",2003,36.1,"Lubelskie"
"Y15-24","PL32",2003,40.5,"Podkarpackie"
"Y15-24","PL33",2003,45.4,"Swietokrzyskie"
"Y15-24","PL34",2003,32.1,"Podlaskie"
"Y15-24","PL4",2003,42.1,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2003,37.9,"Wielkopolskie"
"Y15-24","PL42",2003,48.9,"Zachodniopomorskie"
"Y15-24","PL43",2003,49.7,"Lubuskie"
"Y15-24","PL5",2003,45.1,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2003,45.2,"Dolnoslaskie"
"Y15-24","PL52",2003,44.8,"Opolskie"
"Y15-24","PL6",2003,42.8,"Region Pólnocny"
"Y15-24","PL61",2003,41.7,"Kujawsko-Pomorskie"
"Y15-24","PL62",2003,50.1,"Warminsko-Mazurskie"
"Y15-24","PL63",2003,39.4,"Pomorskie"
"Y15-24","PT",2003,13.5,"Portugal"
"Y15-24","PT1",2003,13.8,"Continente"
"Y15-24","PT11",2003,12.3,"Norte"
"Y15-24","PT15",2003,NA,"Algarve"
"Y15-24","PT16",2003,10.2,"Centro (PT)"
"Y15-24","PT17",2003,17,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2003,20.7,"Alentejo"
"Y15-24","PT2",2003,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2003,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2003,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2003,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2003,19.5,"Romania"
"Y15-24","RO1",2003,19,"Macroregiunea unu"
"Y15-24","RO11",2003,13.7,"Nord-Vest"
"Y15-24","RO12",2003,25.8,"Centru"
"Y15-24","RO2",2003,15.7,"Macroregiunea doi"
"Y15-24","RO21",2003,13.8,"Nord-Est"
"Y15-24","RO22",2003,18.5,"Sud-Est"
"Y15-24","RO3",2003,24.6,"Macroregiunea trei"
"Y15-24","RO31",2003,20.6,"Sud - Muntenia"
"Y15-24","RO32",2003,30.2,"Bucuresti - Ilfov"
"Y15-24","RO4",2003,20.9,"Macroregiunea patru"
"Y15-24","RO41",2003,21,"Sud-Vest Oltenia"
"Y15-24","RO42",2003,20.8,"Vest"
"Y15-24","SE",2003,14.3,"Sweden"
"Y15-24","SE1",2003,14.7,"Östra Sverige"
"Y15-24","SE11",2003,13.8,"Stockholm"
"Y15-24","SE12",2003,15.8,"Östra Mellansverige"
"Y15-24","SE2",2003,13.6,"Södra Sverige"
"Y15-24","SE21",2003,13.3,"Småland med öarna"
"Y15-24","SE22",2003,16.4,"Sydsverige"
"Y15-24","SE23",2003,11.7,"Västsverige"
"Y15-24","SE3",2003,15.3,"Norra Sverige"
"Y15-24","SE31",2003,15.3,"Norra Mellansverige"
"Y15-24","SE32",2003,18.6,"Mellersta Norrland"
"Y15-24","SE33",2003,13.2,"Övre Norrland"
"Y15-24","SI",2003,15.3,"Slovenia"
"Y15-24","SI0",2003,15.3,"Slovenija"
"Y15-24","SI01",2003,19.1,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2003,10.6,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2003,32.9,"Slovakia"
"Y15-24","SK0",2003,32.9,"Slovensko"
"Y15-24","SK01",2003,12.8,"Bratislavský kraj"
"Y15-24","SK02",2003,29.2,"Západné Slovensko"
"Y15-24","SK03",2003,38.1,"Stredné Slovensko"
"Y15-24","SK04",2003,40,"Východné Slovensko"
"Y15-24","UK",2003,11.4,"United Kingdom"
"Y15-24","UKC",2003,16.4,"North East (UK)"
"Y15-24","UKC1",2003,18.6,"Tees Valley and Durham"
"Y15-24","UKC2",2003,14.9,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2003,11.5,"North West (UK)"
"Y15-24","UKD1",2003,NA,"Cumbria"
"Y15-24","UKD3",2003,13.3,"Greater Manchester"
"Y15-24","UKD4",2003,12.1,"Lancashire"
"Y15-24","UKE",2003,12.6,"Yorkshire and The Humber"
"Y15-24","UKE1",2003,NA,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2003,NA,"North Yorkshire"
"Y15-24","UKE3",2003,15.8,"South Yorkshire"
"Y15-24","UKE4",2003,12.5,"West Yorkshire"
"Y15-24","UKF",2003,8.8,"East Midlands (UK)"
"Y15-24","UKF1",2003,8.6,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2003,NA,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2003,NA,"Lincolnshire"
"Y15-24","UKG",2003,13.6,"West Midlands (UK)"
"Y15-24","UKG1",2003,NA,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2003,10.9,"Shropshire and Staffordshire"
"Y15-24","UKG3",2003,17.3,"West Midlands"
"Y15-24","UKH",2003,9.4,"East of England"
"Y15-24","UKH1",2003,8.3,"East Anglia"
"Y15-24","UKH2",2003,NA,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2003,12.2,"Essex"
"Y15-24","UKI",2003,14.3,"London"
"Y15-24","UKI1",2003,16.3,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2003,12.9,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2003,7.6,"South East (UK)"
"Y15-24","UKJ1",2003,7.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2003,8.1,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2003,NA,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2003,NA,"Kent"
"Y15-24","UKK",2003,9.2,"South West (UK)"
"Y15-24","UKK1",2003,8.8,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2003,NA,"Dorset and Somerset"
"Y15-24","UKK3",2003,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2003,NA,"Devon"
"Y15-24","UKL",2003,12.8,"Wales"
"Y15-24","UKL1",2003,13.2,"West Wales and The Valleys"
"Y15-24","UKL2",2003,NA,"East Wales"
"Y15-24","UKM",2003,12.8,"Scotland"
"Y15-24","UKM2",2003,8.5,"Eastern Scotland"
"Y15-24","UKM3",2003,17.6,"South Western Scotland"
"Y15-24","UKM5",2003,NA,"North Eastern Scotland"
"Y15-24","UKM6",2003,NA,"Highlands and Islands"
"Y15-24","UKN",2003,9.9,"Northern Ireland (UK)"
"Y15-24","UKN0",2003,9.9,"Northern Ireland (UK)"
"Y20-64","AT",2003,4.7,"Austria"
"Y20-64","AT1",2003,6,"Ostösterreich"
"Y20-64","AT11",2003,5.7,"Burgenland (AT)"
"Y20-64","AT12",2003,3.8,"Niederösterreich"
"Y20-64","AT13",2003,8.1,"Wien"
"Y20-64","AT2",2003,4,"Südösterreich"
"Y20-64","AT21",2003,4.3,"Kärnten"
"Y20-64","AT22",2003,3.9,"Steiermark"
"Y20-64","AT3",2003,3.5,"Westösterreich"
"Y20-64","AT31",2003,4.1,"Oberösterreich"
"Y20-64","AT32",2003,2.2,"Salzburg"
"Y20-64","AT33",2003,2.9,"Tirol"
"Y20-64","AT34",2003,3.9,"Vorarlberg"
"Y20-64","BE",2003,7.4,"Belgium"
"Y20-64","BE1",2003,14.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2003,14.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2003,4.9,"Vlaams Gewest"
"Y20-64","BE21",2003,6,"Prov. Antwerpen"
"Y20-64","BE22",2003,6.2,"Prov. Limburg (BE)"
"Y20-64","BE23",2003,4.5,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2003,4.2,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2003,3.8,"Prov. West-Vlaanderen"
"Y20-64","BE3",2003,10.2,"Région wallonne"
"Y20-64","BE31",2003,7.3,"Prov. Brabant Wallon"
"Y20-64","BE32",2003,13.2,"Prov. Hainaut"
"Y20-64","BE33",2003,9.8,"Prov. Liège"
"Y20-64","BE34",2003,5.6,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2003,8.4,"Prov. Namur"
"Y20-64","BG",2003,13.6,"Bulgaria"
"Y20-64","BG3",2003,15.6,"Severna i yugoiztochna Bulgaria"
"Y20-64","BG31",2003,11.8,"Severozapaden"
"Y20-64","BG32",2003,14.5,"Severen tsentralen"
"Y20-64","BG33",2003,20.3,"Severoiztochen"
"Y20-64","BG34",2003,15.2,"Yugoiztochen"
"Y20-64","BG4",2003,11.4,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y20-64","BG41",2003,11.2,"Yugozapaden"
"Y20-64","BG42",2003,11.7,"Yuzhen tsentralen"
"Y20-64","CH",2003,4,"Switzerland"
"Y20-64","CH0",2003,4,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2003,5.3,"Région lémanique"
"Y20-64","CH02",2003,3.6,"Espace Mittelland"
"Y20-64","CH03",2003,3.5,"Nordwestschweiz"
"Y20-64","CH04",2003,4.2,"Zürich"
"Y20-64","CH05",2003,3.5,"Ostschweiz"
"Y20-64","CH06",2003,3.7,"Zentralschweiz"
"Y20-64","CH07",2003,4.5,"Ticino"
"Y20-64","CY",2003,4.1,"Cyprus"
"Y20-64","CY0",2003,4.1,"Kypros"
"Y20-64","CY00",2003,4.1,"Kypros"
"Y20-64","CZ",2003,7.3,"Czech Republic"
"Y20-64","CZ0",2003,7.3,"Ceská republika"
"Y20-64","CZ01",2003,4,"Praha"
"Y20-64","CZ02",2003,4.9,"Strední Cechy"
"Y20-64","CZ03",2003,4.7,"Jihozápad"
"Y20-64","CZ04",2003,10.7,"Severozápad"
"Y20-64","CZ05",2003,5.9,"Severovýchod"
"Y20-64","CZ06",2003,6.9,"Jihovýchod"
"Y20-64","CZ07",2003,8.2,"Strední Morava"
"Y20-64","CZ08",2003,13.6,"Moravskoslezsko"
"Y20-64","DE",2003,9.9,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2003,5.8,"Baden-Württemberg"
"Y20-64","DE11",2003,5.9,"Stuttgart"
"Y20-64","DE12",2003,6.2,"Karlsruhe"
"Y20-64","DE13",2003,5.2,"Freiburg"
"Y20-64","DE14",2003,5.5,"Tübingen"
"Y20-64","DE2",2003,6.2,"Bayern"
"Y20-64","DE21",2003,5.1,"Oberbayern"
"Y20-64","DE22",2003,5.7,"Niederbayern"
"Y20-64","DE23",2003,6.7,"Oberpfalz"
"Y20-64","DE24",2003,8.8,"Oberfranken"
"Y20-64","DE25",2003,7.5,"Mittelfranken"
"Y20-64","DE26",2003,6.4,"Unterfranken"
"Y20-64","DE27",2003,5.9,"Schwaben"
"Y20-64","DE3",2003,18.1,"Berlin"
"Y20-64","DE30",2003,18.1,"Berlin"
"Y20-64","DE4",2003,18.7,"Brandenburg"
"Y20-64","DE40",2003,18.7,"Brandenburg"
"Y20-64","DE5",2003,11.4,"Bremen"
"Y20-64","DE50",2003,11.4,"Bremen"
"Y20-64","DE6",2003,9.7,"Hamburg"
"Y20-64","DE60",2003,9.7,"Hamburg"
"Y20-64","DE7",2003,7.1,"Hessen"
"Y20-64","DE71",2003,6.8,"Darmstadt"
"Y20-64","DE72",2003,7.5,"Gießen"
"Y20-64","DE73",2003,7.6,"Kassel"
"Y20-64","DE8",2003,20.9,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2003,20.9,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2003,8.6,"Niedersachsen"
"Y20-64","DE91",2003,10,"Braunschweig"
"Y20-64","DE92",2003,8.3,"Hannover"
"Y20-64","DE93",2003,8.1,"Lüneburg"
"Y20-64","DE94",2003,8.3,"Weser-Ems"
"Y20-64","DEA",2003,8.9,"Nordrhein-Westfalen"
"Y20-64","DEA1",2003,9.1,"Düsseldorf"
"Y20-64","DEA2",2003,7.9,"Köln"
"Y20-64","DEA3",2003,8.7,"Münster"
"Y20-64","DEA4",2003,8.1,"Detmold"
"Y20-64","DEA5",2003,10.1,"Arnsberg"
"Y20-64","DEB",2003,6.3,"Rheinland-Pfalz"
"Y20-64","DEB1",2003,6.6,"Koblenz"
"Y20-64","DEB2",2003,4.8,"Trier"
"Y20-64","DEB3",2003,6.6,"Rheinhessen-Pfalz"
"Y20-64","DEC",2003,8.3,"Saarland"
"Y20-64","DEC0",2003,8.3,"Saarland"
"Y20-64","DED",2003,18.3,"Sachsen"
"Y20-64","DED2",2003,17.1,"Dresden"
"Y20-64","DEE",2003,20.7,"Sachsen-Anhalt"
"Y20-64","DEE0",2003,20.7,"Sachsen-Anhalt"
"Y20-64","DEF",2003,8.6,"Schleswig-Holstein"
"Y20-64","DEF0",2003,8.6,"Schleswig-Holstein"
"Y20-64","DEG",2003,17,"Thüringen"
"Y20-64","DEG0",2003,17,"Thüringen"
"Y20-64","DK",2003,5,"Denmark"
"Y20-64","DK0",2003,5,"Danmark"
"Y20-64","EA17",2003,8.8,"Euro area (17 countries)"
"Y20-64","EA18",2003,8.8,"Euro area (18 countries)"
"Y20-64","EA19",2003,8.8,"Euro area (19 countries)"
"Y20-64","EE",2003,10.9,"Estonia"
"Y20-64","EE0",2003,10.9,"Eesti"
"Y20-64","EE00",2003,10.9,"Eesti"
"Y20-64","EL",2003,9.3,"Greece"
"Y20-64","EL1",2003,10.5,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2003,10,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2003,10,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2003,15.7,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2003,10.3,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2003,9.5,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2003,11,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2003,10,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2003,9.4,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2003,9.7,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2003,8.3,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2003,8.6,"Attiki"
"Y20-64","EL30",2003,8.6,"Attiki"
"Y20-64","EL4",2003,7,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2003,7.5,"Voreio Aigaio"
"Y20-64","EL42",2003,10.7,"Notio Aigaio"
"Y20-64","EL43",2003,4.9,"Kriti"
"Y20-64","ES",2003,10.7,"Spain"
"Y20-64","ES1",2003,11.2,"Noroeste (ES)"
"Y20-64","ES11",2003,11.7,"Galicia"
"Y20-64","ES12",2003,10.6,"Principado de Asturias"
"Y20-64","ES13",2003,9.9,"Cantabria"
"Y20-64","ES2",2003,7.4,"Noreste (ES)"
"Y20-64","ES21",2003,8.9,"País Vasco"
"Y20-64","ES22",2003,5.1,"Comunidad Foral de Navarra"
"Y20-64","ES23",2003,5,"La Rioja"
"Y20-64","ES24",2003,6.3,"Aragón"
"Y20-64","ES3",2003,6.9,"Comunidad de Madrid"
"Y20-64","ES30",2003,6.9,"Comunidad de Madrid"
"Y20-64","ES4",2003,11.5,"Centro (ES)"
"Y20-64","ES41",2003,10.9,"Castilla y León"
"Y20-64","ES42",2003,9.7,"Castilla-la Mancha"
"Y20-64","ES43",2003,16.1,"Extremadura"
"Y20-64","ES5",2003,10,"Este (ES)"
"Y20-64","ES51",2003,9.6,"Cataluña"
"Y20-64","ES52",2003,10.9,"Comunidad Valenciana"
"Y20-64","ES53",2003,8.1,"Illes Balears"
"Y20-64","ES6",2003,15.9,"Sur (ES)"
"Y20-64","ES61",2003,17.3,"Andalucía"
"Y20-64","ES62",2003,8.8,"Región de Murcia"
"Y20-64","ES63",2003,8.4,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2003,NA,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2003,10.7,"Canarias (ES)"
"Y20-64","ES70",2003,10.7,"Canarias (ES)"
"Y20-64","EU15",2003,7.8,"European Union (15 countries)"
"Y20-64","EU27",2003,8.8,"European Union (27 countries)"
"Y20-64","EU28",2003,8.8,"European Union (28 countries)"
"Y20-64","FI",2003,8.8,"Finland"
"Y20-64","FI1",2003,8.8,"Manner-Suomi"
"Y20-64","FI19",2003,8.8,"Länsi-Suomi"
"Y20-64","FI2",2003,NA,"Åland"
"Y20-64","FI20",2003,NA,"Åland"
"Y20-64","FR",2003,8.5,"France"
"Y20-64","FR1",2003,8.1,"Île de France"
"Y20-64","FR10",2003,8.1,"Île de France"
"Y20-64","FR2",2003,7.2,"Bassin Parisien"
"Y20-64","FR21",2003,7.9,"Champagne-Ardenne"
"Y20-64","FR22",2003,9.1,"Picardie"
"Y20-64","FR23",2003,8.5,"Haute-Normandie"
"Y20-64","FR24",2003,5.3,"Centre (FR)"
"Y20-64","FR25",2003,7.5,"Basse-Normandie"
"Y20-64","FR26",2003,6,"Bourgogne"
"Y20-64","FR3",2003,9.8,"Nord - Pas-de-Calais"
"Y20-64","FR30",2003,9.8,"Nord - Pas-de-Calais"
"Y20-64","FR4",2003,7.2,"Est (FR)"
"Y20-64","FR41",2003,8,"Lorraine"
"Y20-64","FR42",2003,6.6,"Alsace"
"Y20-64","FR43",2003,NA,"Franche-Comté"
"Y20-64","FR5",2003,7,"Ouest (FR)"
"Y20-64","FR51",2003,7,"Pays de la Loire"
"Y20-64","FR52",2003,6.6,"Bretagne"
"Y20-64","FR53",2003,7.5,"Poitou-Charentes"
"Y20-64","FR6",2003,8.7,"Sud-Ouest (FR)"
"Y20-64","FR61",2003,8.4,"Aquitaine"
"Y20-64","FR62",2003,9.9,"Midi-Pyrénées"
"Y20-64","FR63",2003,NA,"Limousin"
"Y20-64","FR7",2003,7,"Centre-Est (FR)"
"Y20-64","FR71",2003,7.2,"Rhône-Alpes"
"Y20-64","FR72",2003,NA,"Auvergne"
"Y20-64","FR8",2003,10.5,"Méditerranée"
"Y20-64","FR81",2003,12.2,"Languedoc-Roussillon"
"Y20-64","FR82",2003,9.6,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2003,NA,"Corse"
"Y20-64","FR9",2003,26.3,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2003,25.9,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2003,20.5,"Martinique (NUTS 2010)"
"Y20-64","FR93",2003,23.6,"Guyane (NUTS 2010)"
"Y20-64","FR94",2003,30.3,"Réunion (NUTS 2010)"
"Y20-64","HR",2003,13.5,"Croatia"
"Y20-64","HR0",2003,13.5,"Hrvatska"
"Y20-64","HU",2003,5.6,"Hungary"
"Y20-64","HU1",2003,3.9,"Közép-Magyarország"
"Y20-64","HU10",2003,3.9,"Közép-Magyarország"
"Y20-64","HU2",2003,5.2,"Dunántúl"
"Y20-64","HU21",2003,4.2,"Közép-Dunántúl"
"Y20-64","HU22",2003,4.3,"Nyugat-Dunántúl"
"Y20-64","HU23",2003,7.5,"Dél-Dunántúl"
"Y20-64","HU3",2003,7.2,"Alföld és Észak"
"Y20-64","HU31",2003,9.6,"Észak-Magyarország"
"Y20-64","HU32",2003,6.2,"Észak-Alföld"
"Y20-64","HU33",2003,6.2,"Dél-Alföld"
"Y20-64","IE",2003,4.2,"Ireland"
"Y20-64","IE0",2003,4.2,"Éire/Ireland"
"Y20-64","IE01",2003,5,"Border, Midland and Western"
"Y20-64","IE02",2003,3.9,"Southern and Eastern"
"Y20-64","IS",2003,3.2,"Iceland"
"Y20-64","IS0",2003,3.2,"Ísland"
"Y20-64","IS00",2003,3.2,"Ísland"
"Y20-64","IT",2003,8.5,"Italy"
"Y20-64","ITC",2003,3.9,"Nord-Ovest"
"Y20-64","ITC1",2003,4.4,"Piemonte"
"Y20-64","ITC2",2003,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2003,6.7,"Liguria"
"Y20-64","ITC4",2003,3.2,"Lombardia"
"Y20-64","ITF",2003,16.9,"Sud"
"Y20-64","ITF1",2003,5.6,"Abruzzo"
"Y20-64","ITF2",2003,12.1,"Molise"
"Y20-64","ITF3",2003,20.2,"Campania"
"Y20-64","ITF4",2003,12.7,"Puglia"
"Y20-64","ITF5",2003,16.7,"Basilicata"
"Y20-64","ITF6",2003,24.2,"Calabria"
"Y20-64","ITG",2003,19.4,"Isole"
"Y20-64","ITG1",2003,20.2,"Sicilia"
"Y20-64","ITG2",2003,17,"Sardegna"
"Y20-64","ITH",2003,2.8,"Nord-Est"
"Y20-64","ITH1",2003,1.9,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2003,3.2,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2003,3,"Veneto"
"Y20-64","ITH4",2003,3.6,"Friuli-Venezia Giulia"
"Y20-64","ITI",2003,6.4,"Centro (IT)"
"Y20-64","ITI1",2003,4.5,"Toscana"
"Y20-64","ITI2",2003,5.1,"Umbria"
"Y20-64","ITI4",2003,8.7,"Lazio"
"Y20-64","LT",2003,12.4,"Lithuania"
"Y20-64","LT0",2003,12.4,"Lietuva"
"Y20-64","LT00",2003,12.4,"Lietuva"
"Y20-64","LU",2003,3.6,"Luxembourg"
"Y20-64","LU0",2003,3.6,"Luxembourg"
"Y20-64","LU00",2003,3.6,"Luxembourg"
"Y20-64","LV",2003,11.8,"Latvia"
"Y20-64","LV0",2003,11.8,"Latvija"
"Y20-64","LV00",2003,11.8,"Latvija"
"Y20-64","MT",2003,5.5,"Malta"
"Y20-64","MT0",2003,5.5,"Malta"
"Y20-64","MT00",2003,5.5,"Malta"
"Y20-64","NL",2003,3.2,"Netherlands"
"Y20-64","NL1",2003,3.5,"Noord-Nederland"
"Y20-64","NL11",2003,4.4,"Groningen"
"Y20-64","NL12",2003,3.4,"Friesland (NL)"
"Y20-64","NL13",2003,2.7,"Drenthe"
"Y20-64","NL2",2003,2.8,"Oost-Nederland"
"Y20-64","NL21",2003,3,"Overijssel"
"Y20-64","NL22",2003,2.6,"Gelderland"
"Y20-64","NL23",2003,2.9,"Flevoland"
"Y20-64","NL3",2003,3.3,"West-Nederland"
"Y20-64","NL31",2003,3.5,"Utrecht"
"Y20-64","NL32",2003,3.9,"Noord-Holland"
"Y20-64","NL33",2003,3,"Zuid-Holland"
"Y20-64","NL34",2003,1.8,"Zeeland"
"Y20-64","NL4",2003,3.2,"Zuid-Nederland"
"Y20-64","NL41",2003,2.9,"Noord-Brabant"
"Y20-64","NL42",2003,3.7,"Limburg (NL)"
"Y20-64","NO",2003,3.5,"Norway"
"Y20-64","NO0",2003,3.5,"Norge"
"Y20-64","NO01",2003,3.6,"Oslo og Akershus"
"Y20-64","NO02",2003,3,"Hedmark og Oppland"
"Y20-64","NO03",2003,3.8,"Sør-Østlandet"
"Y20-64","NO04",2003,3.7,"Agder og Rogaland"
"Y20-64","NO05",2003,3.2,"Vestlandet"
"Y20-64","NO06",2003,3.3,"Trøndelag"
"Y20-64","NO07",2003,3.6,"Nord-Norge"
"Y20-64","PL",2003,19.3,"Poland"
"Y20-64","PL1",2003,17.6,"Region Centralny"
"Y20-64","PL11",2003,18.9,"Lódzkie"
"Y20-64","PL12",2003,16.8,"Mazowieckie"
"Y20-64","PL2",2003,18.1,"Region Poludniowy"
"Y20-64","PL21",2003,17.5,"Malopolskie"
"Y20-64","PL22",2003,18.6,"Slaskie"
"Y20-64","PL3",2003,17.2,"Region Wschodni"
"Y20-64","PL31",2003,15.9,"Lubelskie"
"Y20-64","PL32",2003,18.3,"Podkarpackie"
"Y20-64","PL33",2003,17.6,"Swietokrzyskie"
"Y20-64","PL34",2003,17.5,"Podlaskie"
"Y20-64","PL4",2003,19.9,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2003,15.9,"Wielkopolskie"
"Y20-64","PL42",2003,26.3,"Zachodniopomorskie"
"Y20-64","PL43",2003,23.6,"Lubuskie"
"Y20-64","PL5",2003,24,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2003,25.3,"Dolnoslaskie"
"Y20-64","PL52",2003,20,"Opolskie"
"Y20-64","PL6",2003,21.8,"Region Pólnocny"
"Y20-64","PL61",2003,20.9,"Kujawsko-Pomorskie"
"Y20-64","PL62",2003,24.6,"Warminsko-Mazurskie"
"Y20-64","PL63",2003,20.9,"Pomorskie"
"Y20-64","PT",2003,6.2,"Portugal"
"Y20-64","PT1",2003,6.3,"Continente"
"Y20-64","PT11",2003,6.5,"Norte"
"Y20-64","PT15",2003,6.8,"Algarve"
"Y20-64","PT16",2003,3.6,"Centro (PT)"
"Y20-64","PT17",2003,8,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2003,7.3,"Alentejo"
"Y20-64","PT2",2003,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2003,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2003,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2003,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2003,6.8,"Romania"
"Y20-64","RO1",2003,6.2,"Macroregiunea unu"
"Y20-64","RO11",2003,5.5,"Nord-Vest"
"Y20-64","RO12",2003,6.9,"Centru"
"Y20-64","RO2",2003,6.5,"Macroregiunea doi"
"Y20-64","RO21",2003,5.8,"Nord-Est"
"Y20-64","RO22",2003,7.4,"Sud-Est"
"Y20-64","RO3",2003,8.1,"Macroregiunea trei"
"Y20-64","RO31",2003,7.6,"Sud - Muntenia"
"Y20-64","RO32",2003,8.9,"Bucuresti - Ilfov"
"Y20-64","RO4",2003,6.4,"Macroregiunea patru"
"Y20-64","RO41",2003,6.2,"Sud-Vest Oltenia"
"Y20-64","RO42",2003,6.6,"Vest"
"Y20-64","SE",2003,5,"Sweden"
"Y20-64","SE1",2003,4.8,"Östra Sverige"
"Y20-64","SE11",2003,4.6,"Stockholm"
"Y20-64","SE12",2003,5.1,"Östra Mellansverige"
"Y20-64","SE2",2003,4.7,"Södra Sverige"
"Y20-64","SE21",2003,3.6,"Småland med öarna"
"Y20-64","SE22",2003,6.2,"Sydsverige"
"Y20-64","SE23",2003,4.2,"Västsverige"
"Y20-64","SE3",2003,6.2,"Norra Sverige"
"Y20-64","SE31",2003,6.7,"Norra Mellansverige"
"Y20-64","SE32",2003,5.3,"Mellersta Norrland"
"Y20-64","SE33",2003,5.9,"Övre Norrland"
"Y20-64","SI",2003,6.4,"Slovenia"
"Y20-64","SI0",2003,6.4,"Slovenija"
"Y20-64","SI01",2003,7.9,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2003,4.8,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2003,16.3,"Slovakia"
"Y20-64","SK0",2003,16.3,"Slovensko"
"Y20-64","SK01",2003,6.7,"Bratislavský kraj"
"Y20-64","SK02",2003,15,"Západné Slovensko"
"Y20-64","SK03",2003,19.5,"Stredné Slovensko"
"Y20-64","SK04",2003,19.6,"Východné Slovensko"
"Y20-64","UK",2003,4.2,"United Kingdom"
"Y20-64","UKC",2003,5.6,"North East (UK)"
"Y20-64","UKC1",2003,7,"Tees Valley and Durham"
"Y20-64","UKC2",2003,4.6,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2003,4,"North West (UK)"
"Y20-64","UKD1",2003,NA,"Cumbria"
"Y20-64","UKD3",2003,4.3,"Greater Manchester"
"Y20-64","UKD4",2003,2.8,"Lancashire"
"Y20-64","UKE",2003,4.4,"Yorkshire and The Humber"
"Y20-64","UKE1",2003,5.2,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2003,NA,"North Yorkshire"
"Y20-64","UKE3",2003,4.9,"South Yorkshire"
"Y20-64","UKE4",2003,4.6,"West Yorkshire"
"Y20-64","UKF",2003,3.6,"East Midlands (UK)"
"Y20-64","UKF1",2003,4.4,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2003,2.7,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2003,NA,"Lincolnshire"
"Y20-64","UKG",2003,4.7,"West Midlands (UK)"
"Y20-64","UKG1",2003,3.2,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2003,3.2,"Shropshire and Staffordshire"
"Y20-64","UKG3",2003,6.4,"West Midlands"
"Y20-64","UKH",2003,3.3,"East of England"
"Y20-64","UKH1",2003,2.9,"East Anglia"
"Y20-64","UKH2",2003,3.6,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2003,3.5,"Essex"
"Y20-64","UKI",2003,6,"London"
"Y20-64","UKI1",2003,7.9,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2003,4.7,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2003,3.4,"South East (UK)"
"Y20-64","UKJ1",2003,3.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2003,2.6,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2003,3.7,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2003,4.2,"Kent"
"Y20-64","UKK",2003,3.1,"South West (UK)"
"Y20-64","UKK1",2003,3.1,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2003,2.7,"Dorset and Somerset"
"Y20-64","UKK3",2003,NA,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2003,3.2,"Devon"
"Y20-64","UKL",2003,3.5,"Wales"
"Y20-64","UKL1",2003,3.8,"West Wales and The Valleys"
"Y20-64","UKL2",2003,3.1,"East Wales"
"Y20-64","UKM",2003,4.2,"Scotland"
"Y20-64","UKM2",2003,3.4,"Eastern Scotland"
"Y20-64","UKM3",2003,4.8,"South Western Scotland"
"Y20-64","UKM5",2003,NA,"North Eastern Scotland"
"Y20-64","UKM6",2003,5.7,"Highlands and Islands"
"Y20-64","UKN",2003,4.9,"Northern Ireland (UK)"
"Y20-64","UKN0",2003,4.9,"Northern Ireland (UK)"
"Y_GE15","AT",2003,4.8,"Austria"
"Y_GE15","AT1",2003,6.2,"Ostösterreich"
"Y_GE15","AT11",2003,5.8,"Burgenland (AT)"
"Y_GE15","AT12",2003,4,"Niederösterreich"
"Y_GE15","AT13",2003,8.3,"Wien"
"Y_GE15","AT2",2003,4.1,"Südösterreich"
"Y_GE15","AT21",2003,4.3,"Kärnten"
"Y_GE15","AT22",2003,4.1,"Steiermark"
"Y_GE15","AT3",2003,3.5,"Westösterreich"
"Y_GE15","AT31",2003,4,"Oberösterreich"
"Y_GE15","AT32",2003,2.2,"Salzburg"
"Y_GE15","AT33",2003,3.1,"Tirol"
"Y_GE15","AT34",2003,4.3,"Vorarlberg"
"Y_GE15","BE",2003,7.7,"Belgium"
"Y_GE15","BE1",2003,14.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2003,14.7,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2003,5.2,"Vlaams Gewest"
"Y_GE15","BE21",2003,6.1,"Prov. Antwerpen"
"Y_GE15","BE22",2003,6.7,"Prov. Limburg (BE)"
"Y_GE15","BE23",2003,5.1,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2003,4.5,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2003,3.9,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2003,10.3,"Région wallonne"
"Y_GE15","BE31",2003,8.2,"Prov. Brabant Wallon"
"Y_GE15","BE32",2003,13.4,"Prov. Hainaut"
"Y_GE15","BE33",2003,9.6,"Prov. Liège"
"Y_GE15","BE34",2003,5.6,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2003,8.3,"Prov. Namur"
"Y_GE15","BG",2003,13.7,"Bulgaria"
"Y_GE15","BG3",2003,15.8,"Severna i yugoiztochna Bulgaria"
"Y_GE15","BG31",2003,12.1,"Severozapaden"
"Y_GE15","BG32",2003,14.7,"Severen tsentralen"
"Y_GE15","BG33",2003,20.3,"Severoiztochen"
"Y_GE15","BG34",2003,15.4,"Yugoiztochen"
"Y_GE15","BG4",2003,11.5,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE15","BG41",2003,11.3,"Yugozapaden"
"Y_GE15","BG42",2003,11.9,"Yuzhen tsentralen"
"Y_GE15","CH",2003,4.1,"Switzerland"
"Y_GE15","CH0",2003,4.1,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2003,5.5,"Région lémanique"
"Y_GE15","CH02",2003,3.7,"Espace Mittelland"
"Y_GE15","CH03",2003,3.6,"Nordwestschweiz"
"Y_GE15","CH04",2003,4.3,"Zürich"
"Y_GE15","CH05",2003,3.6,"Ostschweiz"
"Y_GE15","CH06",2003,3.8,"Zentralschweiz"
"Y_GE15","CH07",2003,4.5,"Ticino"
"Y_GE15","CY",2003,4.1,"Cyprus"
"Y_GE15","CY0",2003,4.1,"Kypros"
"Y_GE15","CY00",2003,4.1,"Kypros"
"Y_GE15","CZ",2003,7.5,"Czech Republic"
"Y_GE15","CZ0",2003,7.5,"Ceská republika"
"Y_GE15","CZ01",2003,4.2,"Praha"
"Y_GE15","CZ02",2003,5.1,"Strední Cechy"
"Y_GE15","CZ03",2003,5,"Jihozápad"
"Y_GE15","CZ04",2003,11,"Severozápad"
"Y_GE15","CZ05",2003,6.2,"Severovýchod"
"Y_GE15","CZ06",2003,7,"Jihovýchod"
"Y_GE15","CZ07",2003,8.4,"Strední Morava"
"Y_GE15","CZ08",2003,14,"Moravskoslezsko"
"Y_GE15","DE",2003,9.8,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2003,5.7,"Baden-Württemberg"
"Y_GE15","DE11",2003,5.9,"Stuttgart"
"Y_GE15","DE12",2003,6.1,"Karlsruhe"
"Y_GE15","DE13",2003,5.1,"Freiburg"
"Y_GE15","DE14",2003,5.4,"Tübingen"
"Y_GE15","DE2",2003,6.1,"Bayern"
"Y_GE15","DE21",2003,5,"Oberbayern"
"Y_GE15","DE22",2003,5.6,"Niederbayern"
"Y_GE15","DE23",2003,6.4,"Oberpfalz"
"Y_GE15","DE24",2003,8.7,"Oberfranken"
"Y_GE15","DE25",2003,7.4,"Mittelfranken"
"Y_GE15","DE26",2003,6.2,"Unterfranken"
"Y_GE15","DE27",2003,5.8,"Schwaben"
"Y_GE15","DE3",2003,18,"Berlin"
"Y_GE15","DE30",2003,18,"Berlin"
"Y_GE15","DE4",2003,18.3,"Brandenburg"
"Y_GE15","DE40",2003,18.3,"Brandenburg"
"Y_GE15","DE5",2003,11.4,"Bremen"
"Y_GE15","DE50",2003,11.4,"Bremen"
"Y_GE15","DE6",2003,9.6,"Hamburg"
"Y_GE15","DE60",2003,9.6,"Hamburg"
"Y_GE15","DE7",2003,7.1,"Hessen"
"Y_GE15","DE71",2003,6.8,"Darmstadt"
"Y_GE15","DE72",2003,7.5,"Gießen"
"Y_GE15","DE73",2003,7.7,"Kassel"
"Y_GE15","DE8",2003,20.2,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2003,20.2,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2003,8.5,"Niedersachsen"
"Y_GE15","DE91",2003,10,"Braunschweig"
"Y_GE15","DE92",2003,8.1,"Hannover"
"Y_GE15","DE93",2003,8.1,"Lüneburg"
"Y_GE15","DE94",2003,8.1,"Weser-Ems"
"Y_GE15","DEA",2003,8.8,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2003,9.1,"Düsseldorf"
"Y_GE15","DEA2",2003,8,"Köln"
"Y_GE15","DEA3",2003,8.6,"Münster"
"Y_GE15","DEA4",2003,8,"Detmold"
"Y_GE15","DEA5",2003,10,"Arnsberg"
"Y_GE15","DEB",2003,6.3,"Rheinland-Pfalz"
"Y_GE15","DEB1",2003,6.5,"Koblenz"
"Y_GE15","DEB2",2003,4.8,"Trier"
"Y_GE15","DEB3",2003,6.5,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2003,8.3,"Saarland"
"Y_GE15","DEC0",2003,8.3,"Saarland"
"Y_GE15","DED",2003,17.8,"Sachsen"
"Y_GE15","DED2",2003,16.7,"Dresden"
"Y_GE15","DEE",2003,19.9,"Sachsen-Anhalt"
"Y_GE15","DEE0",2003,19.9,"Sachsen-Anhalt"
"Y_GE15","DEF",2003,8.6,"Schleswig-Holstein"
"Y_GE15","DEF0",2003,8.6,"Schleswig-Holstein"
"Y_GE15","DEG",2003,16.3,"Thüringen"
"Y_GE15","DEG0",2003,16.3,"Thüringen"
"Y_GE15","DK",2003,5.4,"Denmark"
"Y_GE15","DK0",2003,5.4,"Danmark"
"Y_GE15","EA17",2003,9,"Euro area (17 countries)"
"Y_GE15","EA18",2003,9,"Euro area (18 countries)"
"Y_GE15","EA19",2003,9,"Euro area (19 countries)"
"Y_GE15","EE",2003,11.3,"Estonia"
"Y_GE15","EE0",2003,11.3,"Eesti"
"Y_GE15","EE00",2003,11.3,"Eesti"
"Y_GE15","EL",2003,9.4,"Greece"
"Y_GE15","EL1",2003,10.6,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2003,10.1,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2003,10,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2003,15.9,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2003,10.4,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2003,9.5,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2003,11.3,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2003,10.3,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2003,9.5,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2003,9.4,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2003,8.2,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2003,8.9,"Attiki"
"Y_GE15","EL30",2003,8.9,"Attiki"
"Y_GE15","EL4",2003,7.4,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2003,7.7,"Voreio Aigaio"
"Y_GE15","EL42",2003,11.2,"Notio Aigaio"
"Y_GE15","EL43",2003,5.3,"Kriti"
"Y_GE15","ES",2003,11.3,"Spain"
"Y_GE15","ES1",2003,11.4,"Noroeste (ES)"
"Y_GE15","ES11",2003,11.9,"Galicia"
"Y_GE15","ES12",2003,10.8,"Principado de Asturias"
"Y_GE15","ES13",2003,10.3,"Cantabria"
"Y_GE15","ES2",2003,7.7,"Noreste (ES)"
"Y_GE15","ES21",2003,9.2,"País Vasco"
"Y_GE15","ES22",2003,5.5,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2003,5.1,"La Rioja"
"Y_GE15","ES24",2003,6.7,"Aragón"
"Y_GE15","ES3",2003,7.1,"Comunidad de Madrid"
"Y_GE15","ES30",2003,7.1,"Comunidad de Madrid"
"Y_GE15","ES4",2003,11.8,"Centro (ES)"
"Y_GE15","ES41",2003,11.2,"Castilla y León"
"Y_GE15","ES42",2003,10.1,"Castilla-la Mancha"
"Y_GE15","ES43",2003,16.5,"Extremadura"
"Y_GE15","ES5",2003,10.8,"Este (ES)"
"Y_GE15","ES51",2003,10.5,"Cataluña"
"Y_GE15","ES52",2003,11.4,"Comunidad Valenciana"
"Y_GE15","ES53",2003,9.4,"Illes Balears"
"Y_GE15","ES6",2003,16.6,"Sur (ES)"
"Y_GE15","ES61",2003,17.9,"Andalucía"
"Y_GE15","ES62",2003,9.8,"Región de Murcia"
"Y_GE15","ES63",2003,9.8,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2003,NA,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2003,11.4,"Canarias (ES)"
"Y_GE15","ES70",2003,11.4,"Canarias (ES)"
"Y_GE15","EU15",2003,8,"European Union (15 countries)"
"Y_GE15","EU27",2003,9,"European Union (27 countries)"
"Y_GE15","EU28",2003,9.1,"European Union (28 countries)"
"Y_GE15","FI",2003,10.5,"Finland"
"Y_GE15","FI1",2003,10.5,"Manner-Suomi"
"Y_GE15","FI19",2003,10.5,"Länsi-Suomi"
"Y_GE15","FI2",2003,NA,"Åland"
"Y_GE15","FI20",2003,NA,"Åland"
"Y_GE15","FR",2003,8.8,"France"
"Y_GE15","FR1",2003,8.4,"Île de France"
"Y_GE15","FR10",2003,8.4,"Île de France"
"Y_GE15","FR2",2003,7.4,"Bassin Parisien"
"Y_GE15","FR21",2003,7.9,"Champagne-Ardenne"
"Y_GE15","FR22",2003,9.3,"Picardie"
"Y_GE15","FR23",2003,8.7,"Haute-Normandie"
"Y_GE15","FR24",2003,5.5,"Centre (FR)"
"Y_GE15","FR25",2003,7.7,"Basse-Normandie"
"Y_GE15","FR26",2003,6.1,"Bourgogne"
"Y_GE15","FR3",2003,10.2,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2003,10.2,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2003,7.9,"Est (FR)"
"Y_GE15","FR41",2003,8.8,"Lorraine"
"Y_GE15","FR42",2003,7.2,"Alsace"
"Y_GE15","FR43",2003,7.5,"Franche-Comté"
"Y_GE15","FR5",2003,7.2,"Ouest (FR)"
"Y_GE15","FR51",2003,7.4,"Pays de la Loire"
"Y_GE15","FR52",2003,6.8,"Bretagne"
"Y_GE15","FR53",2003,7.5,"Poitou-Charentes"
"Y_GE15","FR6",2003,8.9,"Sud-Ouest (FR)"
"Y_GE15","FR61",2003,8.4,"Aquitaine"
"Y_GE15","FR62",2003,10.1,"Midi-Pyrénées"
"Y_GE15","FR63",2003,NA,"Limousin"
"Y_GE15","FR7",2003,7.1,"Centre-Est (FR)"
"Y_GE15","FR71",2003,7.3,"Rhône-Alpes"
"Y_GE15","FR72",2003,NA,"Auvergne"
"Y_GE15","FR8",2003,10.9,"Méditerranée"
"Y_GE15","FR81",2003,12.6,"Languedoc-Roussillon"
"Y_GE15","FR82",2003,10,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2003,NA,"Corse"
"Y_GE15","FR9",2003,27.2,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2003,26.2,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2003,21,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2003,24.3,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2003,31.6,"Réunion (NUTS 2010)"
"Y_GE15","HR",2003,13.9,"Croatia"
"Y_GE15","HR0",2003,13.9,"Hrvatska"
"Y_GE15","HU",2003,5.8,"Hungary"
"Y_GE15","HU1",2003,4.1,"Közép-Magyarország"
"Y_GE15","HU10",2003,4.1,"Közép-Magyarország"
"Y_GE15","HU2",2003,5.4,"Dunántúl"
"Y_GE15","HU21",2003,4.3,"Közép-Dunántúl"
"Y_GE15","HU22",2003,4.6,"Nyugat-Dunántúl"
"Y_GE15","HU23",2003,7.8,"Dél-Dunántúl"
"Y_GE15","HU3",2003,7.5,"Alföld és Észak"
"Y_GE15","HU31",2003,9.8,"Észak-Magyarország"
"Y_GE15","HU32",2003,6.4,"Észak-Alföld"
"Y_GE15","HU33",2003,6.4,"Dél-Alföld"
"Y_GE15","IE",2003,4.5,"Ireland"
"Y_GE15","IE0",2003,4.5,"Éire/Ireland"
"Y_GE15","IE01",2003,5.3,"Border, Midland and Western"
"Y_GE15","IE02",2003,4.2,"Southern and Eastern"
"Y_GE15","IS",2003,4,"Iceland"
"Y_GE15","IS0",2003,4,"Ísland"
"Y_GE15","IS00",2003,4,"Ísland"
"Y_GE15","IT",2003,8.9,"Italy"
"Y_GE15","ITC",2003,4.1,"Nord-Ovest"
"Y_GE15","ITC1",2003,4.8,"Piemonte"
"Y_GE15","ITC2",2003,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2003,6.9,"Liguria"
"Y_GE15","ITC4",2003,3.4,"Lombardia"
"Y_GE15","ITF",2003,17.7,"Sud"
"Y_GE15","ITF1",2003,5.6,"Abruzzo"
"Y_GE15","ITF2",2003,12.6,"Molise"
"Y_GE15","ITF3",2003,21.2,"Campania"
"Y_GE15","ITF4",2003,13.6,"Puglia"
"Y_GE15","ITF5",2003,17,"Basilicata"
"Y_GE15","ITF6",2003,25,"Calabria"
"Y_GE15","ITG",2003,19.8,"Isole"
"Y_GE15","ITG1",2003,20.8,"Sicilia"
"Y_GE15","ITG2",2003,17.3,"Sardegna"
"Y_GE15","ITH",2003,3,"Nord-Est"
"Y_GE15","ITH1",2003,1.8,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2003,3.4,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2003,3.1,"Veneto"
"Y_GE15","ITH4",2003,4,"Friuli-Venezia Giulia"
"Y_GE15","ITI",2003,6.6,"Centro (IT)"
"Y_GE15","ITI1",2003,4.7,"Toscana"
"Y_GE15","ITI2",2003,5.2,"Umbria"
"Y_GE15","ITI4",2003,8.9,"Lazio"
"Y_GE15","LT",2003,12.9,"Lithuania"
"Y_GE15","LT0",2003,12.9,"Lietuva"
"Y_GE15","LT00",2003,12.9,"Lietuva"
"Y_GE15","LU",2003,3.7,"Luxembourg"
"Y_GE15","LU0",2003,3.7,"Luxembourg"
"Y_GE15","LU00",2003,3.7,"Luxembourg"
"Y_GE15","LV",2003,12.1,"Latvia"
"Y_GE15","LV0",2003,12.1,"Latvija"
"Y_GE15","LV00",2003,12.1,"Latvija"
"Y_GE15","MT",2003,7.5,"Malta"
"Y_GE15","MT0",2003,7.5,"Malta"
"Y_GE15","MT00",2003,7.5,"Malta"
"Y_GE15","NL",2003,3.6,"Netherlands"
"Y_GE15","NL1",2003,3.8,"Noord-Nederland"
"Y_GE15","NL11",2003,4.6,"Groningen"
"Y_GE15","NL12",2003,3.5,"Friesland (NL)"
"Y_GE15","NL13",2003,3.2,"Drenthe"
"Y_GE15","NL2",2003,3.3,"Oost-Nederland"
"Y_GE15","NL21",2003,3.2,"Overijssel"
"Y_GE15","NL22",2003,3.2,"Gelderland"
"Y_GE15","NL23",2003,3.6,"Flevoland"
"Y_GE15","NL3",2003,3.7,"West-Nederland"
"Y_GE15","NL31",2003,3.9,"Utrecht"
"Y_GE15","NL32",2003,4.1,"Noord-Holland"
"Y_GE15","NL33",2003,3.5,"Zuid-Holland"
"Y_GE15","NL34",2003,1.9,"Zeeland"
"Y_GE15","NL4",2003,3.6,"Zuid-Nederland"
"Y_GE15","NL41",2003,3.4,"Noord-Brabant"
"Y_GE15","NL42",2003,4,"Limburg (NL)"
"Y_GE15","NO",2003,4.2,"Norway"
"Y_GE15","NO0",2003,4.2,"Norge"
"Y_GE15","NO01",2003,4,"Oslo og Akershus"
"Y_GE15","NO02",2003,3.6,"Hedmark og Oppland"
"Y_GE15","NO03",2003,4.6,"Sør-Østlandet"
"Y_GE15","NO04",2003,4,"Agder og Rogaland"
"Y_GE15","NO05",2003,4.2,"Vestlandet"
"Y_GE15","NO06",2003,4.2,"Trøndelag"
"Y_GE15","NO07",2003,5,"Nord-Norge"
"Y_GE15","PL",2003,19.4,"Poland"
"Y_GE15","PL1",2003,17.5,"Region Centralny"
"Y_GE15","PL11",2003,18.9,"Lódzkie"
"Y_GE15","PL12",2003,16.7,"Mazowieckie"
"Y_GE15","PL2",2003,18.6,"Region Poludniowy"
"Y_GE15","PL21",2003,17.7,"Malopolskie"
"Y_GE15","PL22",2003,19.3,"Slaskie"
"Y_GE15","PL3",2003,17,"Region Wschodni"
"Y_GE15","PL31",2003,15.4,"Lubelskie"
"Y_GE15","PL32",2003,18,"Podkarpackie"
"Y_GE15","PL33",2003,18,"Swietokrzyskie"
"Y_GE15","PL34",2003,17.4,"Podlaskie"
"Y_GE15","PL4",2003,20.2,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2003,16.1,"Wielkopolskie"
"Y_GE15","PL42",2003,26.7,"Zachodniopomorskie"
"Y_GE15","PL43",2003,23.9,"Lubuskie"
"Y_GE15","PL5",2003,24.2,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2003,25.6,"Dolnoslaskie"
"Y_GE15","PL52",2003,20.1,"Opolskie"
"Y_GE15","PL6",2003,22,"Region Pólnocny"
"Y_GE15","PL61",2003,21.3,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2003,25,"Warminsko-Mazurskie"
"Y_GE15","PL63",2003,20.8,"Pomorskie"
"Y_GE15","PT",2003,6.1,"Portugal"
"Y_GE15","PT1",2003,6.3,"Continente"
"Y_GE15","PT11",2003,6.5,"Norte"
"Y_GE15","PT15",2003,6.9,"Algarve"
"Y_GE15","PT16",2003,3.3,"Centro (PT)"
"Y_GE15","PT17",2003,8.3,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2003,7.5,"Alentejo"
"Y_GE15","PT2",2003,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2003,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2003,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2003,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2003,6.9,"Romania"
"Y_GE15","RO1",2003,6.3,"Macroregiunea unu"
"Y_GE15","RO11",2003,5.7,"Nord-Vest"
"Y_GE15","RO12",2003,7,"Centru"
"Y_GE15","RO2",2003,6.5,"Macroregiunea doi"
"Y_GE15","RO21",2003,5.8,"Nord-Est"
"Y_GE15","RO22",2003,7.6,"Sud-Est"
"Y_GE15","RO3",2003,8.3,"Macroregiunea trei"
"Y_GE15","RO31",2003,7.5,"Sud - Muntenia"
"Y_GE15","RO32",2003,9.6,"Bucuresti - Ilfov"
"Y_GE15","RO4",2003,6.7,"Macroregiunea patru"
"Y_GE15","RO41",2003,6.1,"Sud-Vest Oltenia"
"Y_GE15","RO42",2003,7.4,"Vest"
"Y_GE15","SE",2003,5.6,"Sweden"
"Y_GE15","SE1",2003,5.4,"Östra Sverige"
"Y_GE15","SE11",2003,5.1,"Stockholm"
"Y_GE15","SE12",2003,5.7,"Östra Mellansverige"
"Y_GE15","SE2",2003,5.3,"Södra Sverige"
"Y_GE15","SE21",2003,4.2,"Småland med öarna"
"Y_GE15","SE22",2003,6.7,"Sydsverige"
"Y_GE15","SE23",2003,4.8,"Västsverige"
"Y_GE15","SE3",2003,6.5,"Norra Sverige"
"Y_GE15","SE31",2003,6.9,"Norra Mellansverige"
"Y_GE15","SE32",2003,5.9,"Mellersta Norrland"
"Y_GE15","SE33",2003,6.3,"Övre Norrland"
"Y_GE15","SI",2003,6.5,"Slovenia"
"Y_GE15","SI0",2003,6.5,"Slovenija"
"Y_GE15","SI01",2003,7.9,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2003,4.9,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2003,17.1,"Slovakia"
"Y_GE15","SK0",2003,17.1,"Slovensko"
"Y_GE15","SK01",2003,6.9,"Bratislavský kraj"
"Y_GE15","SK02",2003,15.6,"Západné Slovensko"
"Y_GE15","SK03",2003,20.4,"Stredné Slovensko"
"Y_GE15","SK04",2003,20.8,"Východné Slovensko"
"Y_GE15","UK",2003,4.8,"United Kingdom"
"Y_GE15","UKC",2003,6.5,"North East (UK)"
"Y_GE15","UKC1",2003,7.6,"Tees Valley and Durham"
"Y_GE15","UKC2",2003,5.7,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2003,4.7,"North West (UK)"
"Y_GE15","UKD1",2003,4.8,"Cumbria"
"Y_GE15","UKD3",2003,5,"Greater Manchester"
"Y_GE15","UKD4",2003,3.9,"Lancashire"
"Y_GE15","UKE",2003,5.3,"Yorkshire and The Humber"
"Y_GE15","UKE1",2003,6.3,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2003,2.6,"North Yorkshire"
"Y_GE15","UKE3",2003,6.2,"South Yorkshire"
"Y_GE15","UKE4",2003,5.3,"West Yorkshire"
"Y_GE15","UKF",2003,3.9,"East Midlands (UK)"
"Y_GE15","UKF1",2003,4.5,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2003,3.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2003,3.8,"Lincolnshire"
"Y_GE15","UKG",2003,5.5,"West Midlands (UK)"
"Y_GE15","UKG1",2003,3.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2003,4.1,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2003,7.4,"West Midlands"
"Y_GE15","UKH",2003,3.8,"East of England"
"Y_GE15","UKH1",2003,3.5,"East Anglia"
"Y_GE15","UKH2",2003,3.7,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2003,4.4,"Essex"
"Y_GE15","UKI",2003,6.6,"London"
"Y_GE15","UKI1",2003,8.7,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2003,5.3,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2003,3.7,"South East (UK)"
"Y_GE15","UKJ1",2003,3.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2003,2.9,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2003,4,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2003,4.4,"Kent"
"Y_GE15","UKK",2003,3.6,"South West (UK)"
"Y_GE15","UKK1",2003,3.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2003,3.3,"Dorset and Somerset"
"Y_GE15","UKK3",2003,NA,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2003,4,"Devon"
"Y_GE15","UKL",2003,4.4,"Wales"
"Y_GE15","UKL1",2003,4.6,"West Wales and The Valleys"
"Y_GE15","UKL2",2003,3.9,"East Wales"
"Y_GE15","UKM",2003,5.3,"Scotland"
"Y_GE15","UKM2",2003,3.9,"Eastern Scotland"
"Y_GE15","UKM3",2003,6.7,"South Western Scotland"
"Y_GE15","UKM5",2003,NA,"North Eastern Scotland"
"Y_GE15","UKM6",2003,6.5,"Highlands and Islands"
"Y_GE15","UKN",2003,5.2,"Northern Ireland (UK)"
"Y_GE15","UKN0",2003,5.2,"Northern Ireland (UK)"
"Y_GE25","AT",2003,4.4,"Austria"
"Y_GE25","AT1",2003,5.7,"Ostösterreich"
"Y_GE25","AT11",2003,5.3,"Burgenland (AT)"
"Y_GE25","AT12",2003,3.7,"Niederösterreich"
"Y_GE25","AT13",2003,7.6,"Wien"
"Y_GE25","AT2",2003,3.8,"Südösterreich"
"Y_GE25","AT21",2003,3.7,"Kärnten"
"Y_GE25","AT22",2003,3.9,"Steiermark"
"Y_GE25","AT3",2003,3.2,"Westösterreich"
"Y_GE25","AT31",2003,3.6,"Oberösterreich"
"Y_GE25","AT32",2003,2.1,"Salzburg"
"Y_GE25","AT33",2003,2.8,"Tirol"
"Y_GE25","AT34",2003,3.8,"Vorarlberg"
"Y_GE25","BE",2003,6.5,"Belgium"
"Y_GE25","BE1",2003,12.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2003,12.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2003,4.3,"Vlaams Gewest"
"Y_GE25","BE21",2003,5,"Prov. Antwerpen"
"Y_GE25","BE22",2003,5.7,"Prov. Limburg (BE)"
"Y_GE25","BE23",2003,4.2,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2003,3.6,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2003,3.1,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2003,8.8,"Région wallonne"
"Y_GE25","BE31",2003,6.7,"Prov. Brabant Wallon"
"Y_GE25","BE32",2003,11.2,"Prov. Hainaut"
"Y_GE25","BE33",2003,8.5,"Prov. Liège"
"Y_GE25","BE34",2003,NA,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2003,6.7,"Prov. Namur"
"Y_GE25","BG",2003,12.4,"Bulgaria"
"Y_GE25","BG3",2003,14.3,"Severna i yugoiztochna Bulgaria"
"Y_GE25","BG31",2003,10.8,"Severozapaden"
"Y_GE25","BG32",2003,13.1,"Severen tsentralen"
"Y_GE25","BG33",2003,19.1,"Severoiztochen"
"Y_GE25","BG34",2003,13.4,"Yugoiztochen"
"Y_GE25","BG4",2003,10.3,"Yugozapadna i yuzhna tsentralna Bulgaria"
"Y_GE25","BG41",2003,10.3,"Yugozapaden"
"Y_GE25","BG42",2003,10.4,"Yuzhen tsentralen"
"Y_GE25","CH",2003,3.4,"Switzerland"
"Y_GE25","CH0",2003,3.4,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2003,4.4,"Région lémanique"
"Y_GE25","CH02",2003,2.8,"Espace Mittelland"
"Y_GE25","CH03",2003,3,"Nordwestschweiz"
"Y_GE25","CH04",2003,3.8,"Zürich"
"Y_GE25","CH05",2003,2.8,"Ostschweiz"
"Y_GE25","CH06",2003,3.1,"Zentralschweiz"
"Y_GE25","CH07",2003,3.6,"Ticino"
"Y_GE25","CY",2003,3.6,"Cyprus"
"Y_GE25","CY0",2003,3.6,"Kypros"
"Y_GE25","CY00",2003,3.6,"Kypros"
"Y_GE25","CZ",2003,6.5,"Czech Republic"
"Y_GE25","CZ0",2003,6.5,"Ceská republika"
"Y_GE25","CZ01",2003,3.8,"Praha"
"Y_GE25","CZ02",2003,5,"Strední Cechy"
"Y_GE25","CZ03",2003,4.3,"Jihozápad"
"Y_GE25","CZ04",2003,9.9,"Severozápad"
"Y_GE25","CZ05",2003,5.1,"Severovýchod"
"Y_GE25","CZ06",2003,5.7,"Jihovýchod"
"Y_GE25","CZ07",2003,7.1,"Strední Morava"
"Y_GE25","CZ08",2003,12.4,"Moravskoslezsko"
"Y_GE25","DE",2003,9.6,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2003,5.5,"Baden-Württemberg"
"Y_GE25","DE11",2003,5.5,"Stuttgart"
"Y_GE25","DE12",2003,6,"Karlsruhe"
"Y_GE25","DE13",2003,5,"Freiburg"
"Y_GE25","DE14",2003,5.1,"Tübingen"
"Y_GE25","DE2",2003,5.9,"Bayern"
"Y_GE25","DE21",2003,4.9,"Oberbayern"
"Y_GE25","DE22",2003,5.3,"Niederbayern"
"Y_GE25","DE23",2003,6.3,"Oberpfalz"
"Y_GE25","DE24",2003,8.4,"Oberfranken"
"Y_GE25","DE25",2003,7.6,"Mittelfranken"
"Y_GE25","DE26",2003,6,"Unterfranken"
"Y_GE25","DE27",2003,5.6,"Schwaben"
"Y_GE25","DE3",2003,17.6,"Berlin"
"Y_GE25","DE30",2003,17.6,"Berlin"
"Y_GE25","DE4",2003,18.2,"Brandenburg"
"Y_GE25","DE40",2003,18.2,"Brandenburg"
"Y_GE25","DE5",2003,10.7,"Bremen"
"Y_GE25","DE50",2003,10.7,"Bremen"
"Y_GE25","DE6",2003,9.6,"Hamburg"
"Y_GE25","DE60",2003,9.6,"Hamburg"
"Y_GE25","DE7",2003,6.7,"Hessen"
"Y_GE25","DE71",2003,6.5,"Darmstadt"
"Y_GE25","DE72",2003,7,"Gießen"
"Y_GE25","DE73",2003,7.2,"Kassel"
"Y_GE25","DE8",2003,20.3,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2003,20.3,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2003,8.3,"Niedersachsen"
"Y_GE25","DE91",2003,9.6,"Braunschweig"
"Y_GE25","DE92",2003,8.1,"Hannover"
"Y_GE25","DE93",2003,7.8,"Lüneburg"
"Y_GE25","DE94",2003,7.9,"Weser-Ems"
"Y_GE25","DEA",2003,8.6,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2003,8.7,"Düsseldorf"
"Y_GE25","DEA2",2003,7.6,"Köln"
"Y_GE25","DEA3",2003,8.5,"Münster"
"Y_GE25","DEA4",2003,7.8,"Detmold"
"Y_GE25","DEA5",2003,10.2,"Arnsberg"
"Y_GE25","DEB",2003,6.2,"Rheinland-Pfalz"
"Y_GE25","DEB1",2003,6.1,"Koblenz"
"Y_GE25","DEB2",2003,4.9,"Trier"
"Y_GE25","DEB3",2003,6.6,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2003,8,"Saarland"
"Y_GE25","DEC0",2003,8,"Saarland"
"Y_GE25","DED",2003,18,"Sachsen"
"Y_GE25","DED2",2003,16.5,"Dresden"
"Y_GE25","DEE",2003,20.6,"Sachsen-Anhalt"
"Y_GE25","DEE0",2003,20.6,"Sachsen-Anhalt"
"Y_GE25","DEF",2003,8.4,"Schleswig-Holstein"
"Y_GE25","DEF0",2003,8.4,"Schleswig-Holstein"
"Y_GE25","DEG",2003,16.9,"Thüringen"
"Y_GE25","DEG0",2003,16.9,"Thüringen"
"Y_GE25","DK",2003,4.7,"Denmark"
"Y_GE25","DK0",2003,4.7,"Danmark"
"Y_GE25","EA17",2003,7.9,"Euro area (17 countries)"
"Y_GE25","EA18",2003,8,"Euro area (18 countries)"
"Y_GE25","EA19",2003,8,"Euro area (19 countries)"
"Y_GE25","EE",2003,9.3,"Estonia"
"Y_GE25","EE0",2003,9.3,"Eesti"
"Y_GE25","EE00",2003,9.3,"Eesti"
"Y_GE25","EL",2003,7.6,"Greece"
"Y_GE25","EL1",2003,8.8,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2003,8.5,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2003,8.5,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2003,12.8,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2003,8.6,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2003,7.4,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2003,8.6,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2003,7.8,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2003,7,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2003,7.8,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2003,6.6,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2003,7.2,"Attiki"
"Y_GE25","EL30",2003,7.2,"Attiki"
"Y_GE25","EL4",2003,5.4,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2003,5.1,"Voreio Aigaio"
"Y_GE25","EL42",2003,9.5,"Notio Aigaio"
"Y_GE25","EL43",2003,3.4,"Kriti"
"Y_GE25","ES",2003,9.7,"Spain"
"Y_GE25","ES1",2003,10,"Noroeste (ES)"
"Y_GE25","ES11",2003,10.3,"Galicia"
"Y_GE25","ES12",2003,9.4,"Principado de Asturias"
"Y_GE25","ES13",2003,9.2,"Cantabria"
"Y_GE25","ES2",2003,6.6,"Noreste (ES)"
"Y_GE25","ES21",2003,7.8,"País Vasco"
"Y_GE25","ES22",2003,4.5,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2003,4.5,"La Rioja"
"Y_GE25","ES24",2003,5.8,"Aragón"
"Y_GE25","ES3",2003,6.2,"Comunidad de Madrid"
"Y_GE25","ES30",2003,6.2,"Comunidad de Madrid"
"Y_GE25","ES4",2003,10.6,"Centro (ES)"
"Y_GE25","ES41",2003,9.6,"Castilla y León"
"Y_GE25","ES42",2003,9.1,"Castilla-la Mancha"
"Y_GE25","ES43",2003,15.8,"Extremadura"
"Y_GE25","ES5",2003,9,"Este (ES)"
"Y_GE25","ES51",2003,8.6,"Cataluña"
"Y_GE25","ES52",2003,10,"Comunidad Valenciana"
"Y_GE25","ES53",2003,7,"Illes Balears"
"Y_GE25","ES6",2003,14.7,"Sur (ES)"
"Y_GE25","ES61",2003,15.9,"Andalucía"
"Y_GE25","ES62",2003,8.4,"Región de Murcia"
"Y_GE25","ES63",2003,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2003,NA,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2003,9.6,"Canarias (ES)"
"Y_GE25","ES70",2003,9.6,"Canarias (ES)"
"Y_GE25","EU15",2003,7,"European Union (15 countries)"
"Y_GE25","EU27",2003,7.8,"European Union (27 countries)"
"Y_GE25","EU28",2003,7.8,"European Union (28 countries)"
"Y_GE25","FI",2003,7.5,"Finland"
"Y_GE25","FI1",2003,7.6,"Manner-Suomi"
"Y_GE25","FI19",2003,7.5,"Länsi-Suomi"
"Y_GE25","FI2",2003,NA,"Åland"
"Y_GE25","FI20",2003,NA,"Åland"
"Y_GE25","FR",2003,7.7,"France"
"Y_GE25","FR1",2003,7.5,"Île de France"
"Y_GE25","FR10",2003,7.5,"Île de France"
"Y_GE25","FR2",2003,6.5,"Bassin Parisien"
"Y_GE25","FR21",2003,6.8,"Champagne-Ardenne"
"Y_GE25","FR22",2003,8.1,"Picardie"
"Y_GE25","FR23",2003,7.3,"Haute-Normandie"
"Y_GE25","FR24",2003,5,"Centre (FR)"
"Y_GE25","FR25",2003,6.7,"Basse-Normandie"
"Y_GE25","FR26",2003,5.7,"Bourgogne"
"Y_GE25","FR3",2003,8.8,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2003,8.8,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2003,6.2,"Est (FR)"
"Y_GE25","FR41",2003,6.8,"Lorraine"
"Y_GE25","FR42",2003,5.7,"Alsace"
"Y_GE25","FR43",2003,NA,"Franche-Comté"
"Y_GE25","FR5",2003,6.3,"Ouest (FR)"
"Y_GE25","FR51",2003,6.2,"Pays de la Loire"
"Y_GE25","FR52",2003,5.8,"Bretagne"
"Y_GE25","FR53",2003,7.4,"Poitou-Charentes"
"Y_GE25","FR6",2003,7.6,"Sud-Ouest (FR)"
"Y_GE25","FR61",2003,7.5,"Aquitaine"
"Y_GE25","FR62",2003,8.4,"Midi-Pyrénées"
"Y_GE25","FR63",2003,NA,"Limousin"
"Y_GE25","FR7",2003,6.5,"Centre-Est (FR)"
"Y_GE25","FR71",2003,6.7,"Rhône-Alpes"
"Y_GE25","FR72",2003,NA,"Auvergne"
"Y_GE25","FR8",2003,9.7,"Méditerranée"
"Y_GE25","FR81",2003,11.1,"Languedoc-Roussillon"
"Y_GE25","FR82",2003,8.9,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2003,NA,"Corse"
"Y_GE25","FR9",2003,24.1,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2003,23.9,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2003,18.9,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2003,21.5,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2003,27.8,"Réunion (NUTS 2010)"
"Y_GE25","HR",2003,11,"Croatia"
"Y_GE25","HR0",2003,11,"Hrvatska"
"Y_GE25","HU",2003,5,"Hungary"
"Y_GE25","HU1",2003,3.5,"Közép-Magyarország"
"Y_GE25","HU10",2003,3.5,"Közép-Magyarország"
"Y_GE25","HU2",2003,4.7,"Dunántúl"
"Y_GE25","HU21",2003,3.7,"Közép-Dunántúl"
"Y_GE25","HU22",2003,3.8,"Nyugat-Dunántúl"
"Y_GE25","HU23",2003,6.9,"Dél-Dunántúl"
"Y_GE25","HU3",2003,6.5,"Alföld és Észak"
"Y_GE25","HU31",2003,8.6,"Észak-Magyarország"
"Y_GE25","HU32",2003,5.7,"Észak-Alföld"
"Y_GE25","HU33",2003,5.6,"Dél-Alföld"
"Y_GE25","IE",2003,3.7,"Ireland"
"Y_GE25","IE0",2003,3.7,"Éire/Ireland"
"Y_GE25","IE01",2003,4.3,"Border, Midland and Western"
"Y_GE25","IE02",2003,3.5,"Southern and Eastern"
"Y_GE25","IS",2003,2.2,"Iceland"
"Y_GE25","IS0",2003,2.2,"Ísland"
"Y_GE25","IS00",2003,2.2,"Ísland"
"Y_GE25","IT",2003,7.1,"Italy"
"Y_GE25","ITC",2003,3.3,"Nord-Ovest"
"Y_GE25","ITC1",2003,3.8,"Piemonte"
"Y_GE25","ITC2",2003,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2003,5.8,"Liguria"
"Y_GE25","ITC4",2003,2.7,"Lombardia"
"Y_GE25","ITF",2003,14,"Sud"
"Y_GE25","ITF1",2003,5.1,"Abruzzo"
"Y_GE25","ITF2",2003,9.8,"Molise"
"Y_GE25","ITF3",2003,16.3,"Campania"
"Y_GE25","ITF4",2003,10.3,"Puglia"
"Y_GE25","ITF5",2003,14.3,"Basilicata"
"Y_GE25","ITF6",2003,21.3,"Calabria"
"Y_GE25","ITG",2003,16.1,"Isole"
"Y_GE25","ITG1",2003,16.8,"Sicilia"
"Y_GE25","ITG2",2003,14.2,"Sardegna"
"Y_GE25","ITH",2003,2.6,"Nord-Est"
"Y_GE25","ITH1",2003,1.8,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2003,2.9,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2003,2.7,"Veneto"
"Y_GE25","ITH4",2003,3.2,"Friuli-Venezia Giulia"
"Y_GE25","ITI",2003,5.2,"Centro (IT)"
"Y_GE25","ITI1",2003,3.9,"Toscana"
"Y_GE25","ITI2",2003,4.1,"Umbria"
"Y_GE25","ITI4",2003,6.9,"Lazio"
"Y_GE25","LT",2003,11.4,"Lithuania"
"Y_GE25","LT0",2003,11.4,"Lietuva"
"Y_GE25","LT00",2003,11.4,"Lietuva"
"Y_GE25","LU",2003,3.1,"Luxembourg"
"Y_GE25","LU0",2003,3.1,"Luxembourg"
"Y_GE25","LU00",2003,3.1,"Luxembourg"
"Y_GE25","LV",2003,10.9,"Latvia"
"Y_GE25","LV0",2003,10.9,"Latvija"
"Y_GE25","LV00",2003,10.9,"Latvija"
"Y_GE25","MT",2003,4.6,"Malta"
"Y_GE25","MT0",2003,4.6,"Malta"
"Y_GE25","MT00",2003,4.6,"Malta"
"Y_GE25","NL",2003,3,"Netherlands"
"Y_GE25","NL1",2003,3.2,"Noord-Nederland"
"Y_GE25","NL11",2003,4,"Groningen"
"Y_GE25","NL12",2003,3,"Friesland (NL)"
"Y_GE25","NL13",2003,2.5,"Drenthe"
"Y_GE25","NL2",2003,2.6,"Oost-Nederland"
"Y_GE25","NL21",2003,2.7,"Overijssel"
"Y_GE25","NL22",2003,2.6,"Gelderland"
"Y_GE25","NL23",2003,3,"Flevoland"
"Y_GE25","NL3",2003,3.1,"West-Nederland"
"Y_GE25","NL31",2003,3.3,"Utrecht"
"Y_GE25","NL32",2003,3.4,"Noord-Holland"
"Y_GE25","NL33",2003,2.8,"Zuid-Holland"
"Y_GE25","NL34",2003,1.9,"Zeeland"
"Y_GE25","NL4",2003,3.1,"Zuid-Nederland"
"Y_GE25","NL41",2003,2.8,"Noord-Brabant"
"Y_GE25","NL42",2003,3.6,"Limburg (NL)"
"Y_GE25","NO",2003,3,"Norway"
"Y_GE25","NO0",2003,3,"Norge"
"Y_GE25","NO01",2003,3.3,"Oslo og Akershus"
"Y_GE25","NO02",2003,2.5,"Hedmark og Oppland"
"Y_GE25","NO03",2003,3,"Sør-Østlandet"
"Y_GE25","NO04",2003,3.1,"Agder og Rogaland"
"Y_GE25","NO05",2003,2.5,"Vestlandet"
"Y_GE25","NO06",2003,3.2,"Trøndelag"
"Y_GE25","NO07",2003,3,"Nord-Norge"
"Y_GE25","PL",2003,16.1,"Poland"
"Y_GE25","PL1",2003,14.5,"Region Centralny"
"Y_GE25","PL11",2003,15.8,"Lódzkie"
"Y_GE25","PL12",2003,13.8,"Mazowieckie"
"Y_GE25","PL2",2003,14.6,"Region Poludniowy"
"Y_GE25","PL21",2003,13.9,"Malopolskie"
"Y_GE25","PL22",2003,15.2,"Slaskie"
"Y_GE25","PL3",2003,14.1,"Region Wschodni"
"Y_GE25","PL31",2003,12.2,"Lubelskie"
"Y_GE25","PL32",2003,15.2,"Podkarpackie"
"Y_GE25","PL33",2003,14.9,"Swietokrzyskie"
"Y_GE25","PL34",2003,15.3,"Podlaskie"
"Y_GE25","PL4",2003,16.7,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2003,12.2,"Wielkopolskie"
"Y_GE25","PL42",2003,23.8,"Zachodniopomorskie"
"Y_GE25","PL43",2003,20.2,"Lubuskie"
"Y_GE25","PL5",2003,21.1,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2003,22.5,"Dolnoslaskie"
"Y_GE25","PL52",2003,16.8,"Opolskie"
"Y_GE25","PL6",2003,18.9,"Region Pólnocny"
"Y_GE25","PL61",2003,18.3,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2003,21.3,"Warminsko-Mazurskie"
"Y_GE25","PL63",2003,18.1,"Pomorskie"
"Y_GE25","PT",2003,5.2,"Portugal"
"Y_GE25","PT1",2003,5.3,"Continente"
"Y_GE25","PT11",2003,5.6,"Norte"
"Y_GE25","PT15",2003,5.7,"Algarve"
"Y_GE25","PT16",2003,2.7,"Centro (PT)"
"Y_GE25","PT17",2003,7.3,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2003,6,"Alentejo"
"Y_GE25","PT2",2003,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2003,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2003,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2003,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2003,5.4,"Romania"
"Y_GE25","RO1",2003,4.6,"Macroregiunea unu"
"Y_GE25","RO11",2003,4.5,"Nord-Vest"
"Y_GE25","RO12",2003,4.7,"Centru"
"Y_GE25","RO2",2003,5.2,"Macroregiunea doi"
"Y_GE25","RO21",2003,4.6,"Nord-Est"
"Y_GE25","RO22",2003,6.2,"Sud-Est"
"Y_GE25","RO3",2003,6.4,"Macroregiunea trei"
"Y_GE25","RO31",2003,6.1,"Sud - Muntenia"
"Y_GE25","RO32",2003,7,"Bucuresti - Ilfov"
"Y_GE25","RO4",2003,5.1,"Macroregiunea patru"
"Y_GE25","RO41",2003,4.3,"Sud-Vest Oltenia"
"Y_GE25","RO42",2003,6.1,"Vest"
"Y_GE25","SE",2003,4.4,"Sweden"
"Y_GE25","SE1",2003,4.2,"Östra Sverige"
"Y_GE25","SE11",2003,4.1,"Stockholm"
"Y_GE25","SE12",2003,4.3,"Östra Mellansverige"
"Y_GE25","SE2",2003,4.2,"Södra Sverige"
"Y_GE25","SE21",2003,3,"Småland med öarna"
"Y_GE25","SE22",2003,5.4,"Sydsverige"
"Y_GE25","SE23",2003,3.9,"Västsverige"
"Y_GE25","SE3",2003,5.3,"Norra Sverige"
"Y_GE25","SE31",2003,5.8,"Norra Mellansverige"
"Y_GE25","SE32",2003,4.4,"Mellersta Norrland"
"Y_GE25","SE33",2003,5.4,"Övre Norrland"
"Y_GE25","SI",2003,5.5,"Slovenia"
"Y_GE25","SI0",2003,5.5,"Slovenija"
"Y_GE25","SI01",2003,6.6,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2003,4.2,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2003,14.5,"Slovakia"
"Y_GE25","SK0",2003,14.5,"Slovensko"
"Y_GE25","SK01",2003,6,"Bratislavský kraj"
"Y_GE25","SK02",2003,13.5,"Západné Slovensko"
"Y_GE25","SK03",2003,17.4,"Stredné Slovensko"
"Y_GE25","SK04",2003,17.4,"Východné Slovensko"
"Y_GE25","UK",2003,3.7,"United Kingdom"
"Y_GE25","UKC",2003,4.6,"North East (UK)"
"Y_GE25","UKC1",2003,5.7,"Tees Valley and Durham"
"Y_GE25","UKC2",2003,3.9,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2003,3.5,"North West (UK)"
"Y_GE25","UKD1",2003,NA,"Cumbria"
"Y_GE25","UKD3",2003,3.4,"Greater Manchester"
"Y_GE25","UKD4",2003,2.4,"Lancashire"
"Y_GE25","UKE",2003,3.8,"Yorkshire and The Humber"
"Y_GE25","UKE1",2003,5.1,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2003,NA,"North Yorkshire"
"Y_GE25","UKE3",2003,3.9,"South Yorkshire"
"Y_GE25","UKE4",2003,4,"West Yorkshire"
"Y_GE25","UKF",2003,3.1,"East Midlands (UK)"
"Y_GE25","UKF1",2003,3.8,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2003,2.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2003,NA,"Lincolnshire"
"Y_GE25","UKG",2003,4,"West Midlands (UK)"
"Y_GE25","UKG1",2003,3,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2003,2.9,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2003,5.3,"West Midlands"
"Y_GE25","UKH",2003,2.9,"East of England"
"Y_GE25","UKH1",2003,2.7,"East Anglia"
"Y_GE25","UKH2",2003,3.1,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2003,3.1,"Essex"
"Y_GE25","UKI",2003,5.4,"London"
"Y_GE25","UKI1",2003,7.4,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2003,4.1,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2003,3,"South East (UK)"
"Y_GE25","UKJ1",2003,3.1,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2003,2.1,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2003,3.4,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2003,4,"Kent"
"Y_GE25","UKK",2003,2.6,"South West (UK)"
"Y_GE25","UKK1",2003,2.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2003,2.3,"Dorset and Somerset"
"Y_GE25","UKK3",2003,NA,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2003,2.8,"Devon"
"Y_GE25","UKL",2003,2.8,"Wales"
"Y_GE25","UKL1",2003,3,"West Wales and The Valleys"
"Y_GE25","UKL2",2003,2.5,"East Wales"
"Y_GE25","UKM",2003,4,"Scotland"
"Y_GE25","UKM2",2003,3.1,"Eastern Scotland"
"Y_GE25","UKM3",2003,4.4,"South Western Scotland"
"Y_GE25","UKM5",2003,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2003,5.8,"Highlands and Islands"
"Y_GE25","UKN",2003,4.2,"Northern Ireland (UK)"
"Y_GE25","UKN0",2003,4.2,"Northern Ireland (UK)"
"Y15-24","AT",2002,7.2,"Austria"
"Y15-24","AT1",2002,9,"Ostösterreich"
"Y15-24","AT11",2002,NA,"Burgenland (AT)"
"Y15-24","AT12",2002,6.8,"Niederösterreich"
"Y15-24","AT13",2002,11.7,"Wien"
"Y15-24","AT2",2002,7.9,"Südösterreich"
"Y15-24","AT21",2002,NA,"Kärnten"
"Y15-24","AT22",2002,7.4,"Steiermark"
"Y15-24","AT3",2002,5.1,"Westösterreich"
"Y15-24","AT31",2002,5.4,"Oberösterreich"
"Y15-24","AT32",2002,NA,"Salzburg"
"Y15-24","AT33",2002,NA,"Tirol"
"Y15-24","AT34",2002,NA,"Vorarlberg"
"Y15-24","BE",2002,15.7,"Belgium"
"Y15-24","BE1",2002,30.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2002,30.5,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2002,10.6,"Vlaams Gewest"
"Y15-24","BE21",2002,9.9,"Prov. Antwerpen"
"Y15-24","BE22",2002,NA,"Prov. Limburg (BE)"
"Y15-24","BE23",2002,14.8,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2002,12.5,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2002,NA,"Prov. West-Vlaanderen"
"Y15-24","BE3",2002,22.4,"Région wallonne"
"Y15-24","BE31",2002,NA,"Prov. Brabant Wallon"
"Y15-24","BE32",2002,28.3,"Prov. Hainaut"
"Y15-24","BE33",2002,17.2,"Prov. Liège"
"Y15-24","BE34",2002,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2002,NA,"Prov. Namur"
"Y15-24","BG",2002,35.6,"Bulgaria"
"Y15-24","BG41",2002,26.9,"Yugozapaden"
"Y15-24","CH",2002,5.6,"Switzerland"
"Y15-24","CH0",2002,5.6,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2002,7.6,"Région lémanique"
"Y15-24","CH02",2002,4.7,"Espace Mittelland"
"Y15-24","CH03",2002,3.4,"Nordwestschweiz"
"Y15-24","CH04",2002,7.2,"Zürich"
"Y15-24","CH05",2002,6.6,"Ostschweiz"
"Y15-24","CH06",2002,NA,"Zentralschweiz"
"Y15-24","CH07",2002,NA,"Ticino"
"Y15-24","CY",2002,7.7,"Cyprus"
"Y15-24","CY0",2002,7.7,"Kypros"
"Y15-24","CY00",2002,7.7,"Kypros"
"Y15-24","CZ",2002,15.4,"Czech Republic"
"Y15-24","CZ0",2002,15.4,"Ceská republika"
"Y15-24","CZ01",2002,9.1,"Praha"
"Y15-24","CZ02",2002,8,"Strední Cechy"
"Y15-24","CZ03",2002,8,"Jihozápad"
"Y15-24","CZ04",2002,26.3,"Severozápad"
"Y15-24","CZ05",2002,10,"Severovýchod"
"Y15-24","CZ06",2002,15.3,"Jihovýchod"
"Y15-24","CZ07",2002,19.8,"Strední Morava"
"Y15-24","CZ08",2002,25.6,"Moravskoslezsko"
"Y15-24","DE",2002,9.3,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2002,5.4,"Baden-Württemberg"
"Y15-24","DE11",2002,5.3,"Stuttgart"
"Y15-24","DE12",2002,6.8,"Karlsruhe"
"Y15-24","DE13",2002,5.3,"Freiburg"
"Y15-24","DE14",2002,NA,"Tübingen"
"Y15-24","DE2",2002,5.2,"Bayern"
"Y15-24","DE21",2002,3.6,"Oberbayern"
"Y15-24","DE22",2002,6,"Niederbayern"
"Y15-24","DE23",2002,NA,"Oberpfalz"
"Y15-24","DE24",2002,NA,"Oberfranken"
"Y15-24","DE25",2002,5.8,"Mittelfranken"
"Y15-24","DE26",2002,6.6,"Unterfranken"
"Y15-24","DE27",2002,4.6,"Schwaben"
"Y15-24","DE3",2002,19.4,"Berlin"
"Y15-24","DE30",2002,19.4,"Berlin"
"Y15-24","DE4",2002,16.4,"Brandenburg"
"Y15-24","DE40",2002,16.4,"Brandenburg"
"Y15-24","DE5",2002,NA,"Bremen"
"Y15-24","DE50",2002,NA,"Bremen"
"Y15-24","DE6",2002,9.9,"Hamburg"
"Y15-24","DE60",2002,9.9,"Hamburg"
"Y15-24","DE7",2002,7.5,"Hessen"
"Y15-24","DE71",2002,7,"Darmstadt"
"Y15-24","DE72",2002,NA,"Gießen"
"Y15-24","DE73",2002,9.4,"Kassel"
"Y15-24","DE8",2002,14.7,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2002,14.7,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2002,9.1,"Niedersachsen"
"Y15-24","DE91",2002,9.9,"Braunschweig"
"Y15-24","DE92",2002,9.4,"Hannover"
"Y15-24","DE93",2002,10.4,"Lüneburg"
"Y15-24","DE94",2002,7.6,"Weser-Ems"
"Y15-24","DEA",2002,8.4,"Nordrhein-Westfalen"
"Y15-24","DEA1",2002,8.3,"Düsseldorf"
"Y15-24","DEA2",2002,7,"Köln"
"Y15-24","DEA3",2002,8.4,"Münster"
"Y15-24","DEA4",2002,10.6,"Detmold"
"Y15-24","DEA5",2002,8.7,"Arnsberg"
"Y15-24","DEB",2002,7.7,"Rheinland-Pfalz"
"Y15-24","DEB1",2002,7.6,"Koblenz"
"Y15-24","DEB2",2002,NA,"Trier"
"Y15-24","DEB3",2002,8.8,"Rheinhessen-Pfalz"
"Y15-24","DEC",2002,10.7,"Saarland"
"Y15-24","DEC0",2002,10.7,"Saarland"
"Y15-24","DED",2002,14.5,"Sachsen"
"Y15-24","DED2",2002,16.8,"Dresden"
"Y15-24","DEE",2002,14.9,"Sachsen-Anhalt"
"Y15-24","DEE0",2002,14.9,"Sachsen-Anhalt"
"Y15-24","DEF",2002,10.7,"Schleswig-Holstein"
"Y15-24","DEF0",2002,10.7,"Schleswig-Holstein"
"Y15-24","DEG",2002,11.3,"Thüringen"
"Y15-24","DEG0",2002,11.3,"Thüringen"
"Y15-24","DK",2002,7.1,"Denmark"
"Y15-24","DK0",2002,7.1,"Danmark"
"Y15-24","EA17",2002,16.6,"Euro area (17 countries)"
"Y15-24","EA18",2002,16.7,"Euro area (18 countries)"
"Y15-24","EA19",2002,16.7,"Euro area (19 countries)"
"Y15-24","EE",2002,20.2,"Estonia"
"Y15-24","EE0",2002,20.2,"Eesti"
"Y15-24","EE00",2002,20.2,"Eesti"
"Y15-24","EL",2002,25.8,"Greece"
"Y15-24","EL1",2002,28,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2002,24.3,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2002,26.8,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2002,35.2,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2002,32.8,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2002,28.7,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2002,37.4,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2002,NA,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2002,29.5,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2002,29.4,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2002,26.5,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2002,22,"Attiki"
"Y15-24","EL30",2002,22,"Attiki"
"Y15-24","EL4",2002,28.4,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2002,30.6,"Voreio Aigaio"
"Y15-24","EL42",2002,33.8,"Notio Aigaio"
"Y15-24","EL43",2002,24,"Kriti"
"Y15-24","ES",2002,21.5,"Spain"
"Y15-24","ES1",2002,24.1,"Noroeste (ES)"
"Y15-24","ES11",2002,24.9,"Galicia"
"Y15-24","ES12",2002,23,"Principado de Asturias"
"Y15-24","ES13",2002,22,"Cantabria"
"Y15-24","ES2",2002,16.4,"Noreste (ES)"
"Y15-24","ES21",2002,20.6,"País Vasco"
"Y15-24","ES22",2002,12.4,"Comunidad Foral de Navarra"
"Y15-24","ES23",2002,14.5,"La Rioja"
"Y15-24","ES24",2002,12.1,"Aragón"
"Y15-24","ES3",2002,14.3,"Comunidad de Madrid"
"Y15-24","ES30",2002,14.3,"Comunidad de Madrid"
"Y15-24","ES4",2002,22.5,"Centro (ES)"
"Y15-24","ES41",2002,24.7,"Castilla y León"
"Y15-24","ES42",2002,17.6,"Castilla-la Mancha"
"Y15-24","ES43",2002,27.6,"Extremadura"
"Y15-24","ES5",2002,19.9,"Este (ES)"
"Y15-24","ES51",2002,19.7,"Cataluña"
"Y15-24","ES52",2002,21.3,"Comunidad Valenciana"
"Y15-24","ES53",2002,14.5,"Illes Balears"
"Y15-24","ES6",2002,27.7,"Sur (ES)"
"Y15-24","ES61",2002,29.4,"Andalucía"
"Y15-24","ES62",2002,20.2,"Región de Murcia"
"Y15-24","ES63",2002,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES7",2002,20.7,"Canarias (ES)"
"Y15-24","ES70",2002,20.7,"Canarias (ES)"
"Y15-24","EU15",2002,14.8,"European Union (15 countries)"
"Y15-24","EU27",2002,18,"European Union (27 countries)"
"Y15-24","EU28",2002,18.2,"European Union (28 countries)"
"Y15-24","FI",2002,28.2,"Finland"
"Y15-24","FI1",2002,28.2,"Manner-Suomi"
"Y15-24","FI19",2002,29.6,"Länsi-Suomi"
"Y15-24","FI2",2002,NA,"Åland"
"Y15-24","FI20",2002,NA,"Åland"
"Y15-24","FR",2002,19.8,"France"
"Y15-24","FR1",2002,15,"Île de France"
"Y15-24","FR10",2002,15,"Île de France"
"Y15-24","FR2",2002,19.6,"Bassin Parisien"
"Y15-24","FR21",2002,27,"Champagne-Ardenne"
"Y15-24","FR22",2002,20.6,"Picardie"
"Y15-24","FR23",2002,22.2,"Haute-Normandie"
"Y15-24","FR24",2002,16,"Centre (FR)"
"Y15-24","FR25",2002,NA,"Basse-Normandie"
"Y15-24","FR26",2002,NA,"Bourgogne"
"Y15-24","FR3",2002,29.4,"Nord - Pas-de-Calais"
"Y15-24","FR30",2002,29.4,"Nord - Pas-de-Calais"
"Y15-24","FR4",2002,18,"Est (FR)"
"Y15-24","FR41",2002,19.9,"Lorraine"
"Y15-24","FR42",2002,13.4,"Alsace"
"Y15-24","FR43",2002,21.8,"Franche-Comté"
"Y15-24","FR5",2002,15.6,"Ouest (FR)"
"Y15-24","FR51",2002,14.6,"Pays de la Loire"
"Y15-24","FR52",2002,16,"Bretagne"
"Y15-24","FR53",2002,17,"Poitou-Charentes"
"Y15-24","FR6",2002,18.3,"Sud-Ouest (FR)"
"Y15-24","FR61",2002,18.8,"Aquitaine"
"Y15-24","FR62",2002,17.6,"Midi-Pyrénées"
"Y15-24","FR63",2002,NA,"Limousin"
"Y15-24","FR7",2002,16.5,"Centre-Est (FR)"
"Y15-24","FR71",2002,17,"Rhône-Alpes"
"Y15-24","FR72",2002,NA,"Auvergne"
"Y15-24","FR8",2002,24.9,"Méditerranée"
"Y15-24","FR81",2002,31.3,"Languedoc-Roussillon"
"Y15-24","FR82",2002,21.4,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2002,NA,"Corse"
"Y15-24","FR9",2002,51.3,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2002,57.8,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2002,55.2,"Martinique (NUTS 2010)"
"Y15-24","FR93",2002,46.5,"Guyane (NUTS 2010)"
"Y15-24","FR94",2002,48.6,"Réunion (NUTS 2010)"
"Y15-24","HR",2002,36.3,"Croatia"
"Y15-24","HR0",2002,36.3,"Hrvatska"
"Y15-24","HU",2002,11.4,"Hungary"
"Y15-24","HU1",2002,7.9,"Közép-Magyarország"
"Y15-24","HU10",2002,7.9,"Közép-Magyarország"
"Y15-24","HU2",2002,11.5,"Dunántúl"
"Y15-24","HU21",2002,10.7,"Közép-Dunántúl"
"Y15-24","HU22",2002,8.4,"Nyugat-Dunántúl"
"Y15-24","HU23",2002,16.6,"Dél-Dunántúl"
"Y15-24","HU3",2002,13.8,"Alföld és Észak"
"Y15-24","HU31",2002,17.6,"Észak-Magyarország"
"Y15-24","HU32",2002,12.9,"Észak-Alföld"
"Y15-24","HU33",2002,11.5,"Dél-Alföld"
"Y15-24","IE",2002,7.8,"Ireland"
"Y15-24","IE0",2002,7.8,"Éire/Ireland"
"Y15-24","IE01",2002,10.2,"Border, Midland and Western"
"Y15-24","IE02",2002,7.1,"Southern and Eastern"
"Y15-24","IS",2002,6.4,"Iceland"
"Y15-24","IS0",2002,6.4,"Ísland"
"Y15-24","IS00",2002,6.4,"Ísland"
"Y15-24","IT",2002,27.1,"Italy"
"Y15-24","ITC",2002,13.9,"Nord-Ovest"
"Y15-24","ITC1",2002,16.9,"Piemonte"
"Y15-24","ITC2",2002,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2002,24,"Liguria"
"Y15-24","ITC4",2002,11.6,"Lombardia"
"Y15-24","ITF",2002,48.1,"Sud"
"Y15-24","ITF1",2002,17.1,"Abruzzo"
"Y15-24","ITF2",2002,33.4,"Molise"
"Y15-24","ITF3",2002,58.5,"Campania"
"Y15-24","ITF4",2002,36.9,"Puglia"
"Y15-24","ITF5",2002,42.5,"Basilicata"
"Y15-24","ITF6",2002,58.3,"Calabria"
"Y15-24","ITG",2002,49.2,"Isole"
"Y15-24","ITG1",2002,49.7,"Sicilia"
"Y15-24","ITG2",2002,47.9,"Sardegna"
"Y15-24","ITH",2002,7.3,"Nord-Est"
"Y15-24","ITH1",2002,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2002,NA,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2002,7,"Veneto"
"Y15-24","ITH4",2002,9.3,"Friuli-Venezia Giulia"
"Y15-24","ITI",2002,22.6,"Centro (IT)"
"Y15-24","ITI1",2002,17,"Toscana"
"Y15-24","ITI2",2002,15.2,"Umbria"
"Y15-24","ITI4",2002,33.1,"Lazio"
"Y15-24","LT",2002,20.4,"Lithuania"
"Y15-24","LT0",2002,20.4,"Lietuva"
"Y15-24","LT00",2002,20.4,"Lietuva"
"Y15-24","LU",2002,7,"Luxembourg"
"Y15-24","LU0",2002,7,"Luxembourg"
"Y15-24","LU00",2002,7,"Luxembourg"
"Y15-24","LV",2002,25.3,"Latvia"
"Y15-24","LV0",2002,25.3,"Latvija"
"Y15-24","LV00",2002,25.3,"Latvija"
"Y15-24","MT",2002,15.3,"Malta"
"Y15-24","MT0",2002,15.3,"Malta"
"Y15-24","MT00",2002,15.3,"Malta"
"Y15-24","NL",2002,4.6,"Netherlands"
"Y15-24","NL1",2002,6.1,"Noord-Nederland"
"Y15-24","NL11",2002,6.5,"Groningen"
"Y15-24","NL12",2002,5,"Friesland (NL)"
"Y15-24","NL13",2002,7.2,"Drenthe"
"Y15-24","NL2",2002,4.5,"Oost-Nederland"
"Y15-24","NL21",2002,4.3,"Overijssel"
"Y15-24","NL22",2002,4.1,"Gelderland"
"Y15-24","NL23",2002,7,"Flevoland"
"Y15-24","NL3",2002,4,"West-Nederland"
"Y15-24","NL31",2002,4.2,"Utrecht"
"Y15-24","NL32",2002,4.2,"Noord-Holland"
"Y15-24","NL33",2002,3.9,"Zuid-Holland"
"Y15-24","NL34",2002,NA,"Zeeland"
"Y15-24","NL4",2002,5.1,"Zuid-Nederland"
"Y15-24","NL41",2002,4.8,"Noord-Brabant"
"Y15-24","NL42",2002,5.8,"Limburg (NL)"
"Y15-24","NO",2002,13,"Norway"
"Y15-24","NO0",2002,13,"Norge"
"Y15-24","NO01",2002,11,"Oslo og Akershus"
"Y15-24","NO02",2002,15.2,"Hedmark og Oppland"
"Y15-24","NO03",2002,12.3,"Sør-Østlandet"
"Y15-24","NO04",2002,11.8,"Agder og Rogaland"
"Y15-24","NO05",2002,12.1,"Vestlandet"
"Y15-24","NO06",2002,18,"Trøndelag"
"Y15-24","NO07",2002,16.5,"Nord-Norge"
"Y15-24","PL",2002,41.6,"Poland"
"Y15-24","PL1",2002,35.1,"Region Centralny"
"Y15-24","PL11",2002,41.9,"Lódzkie"
"Y15-24","PL12",2002,31.2,"Mazowieckie"
"Y15-24","PL2",2002,39.8,"Region Poludniowy"
"Y15-24","PL21",2002,35.2,"Malopolskie"
"Y15-24","PL22",2002,43.8,"Slaskie"
"Y15-24","PL3",2002,39.7,"Region Wschodni"
"Y15-24","PL31",2002,36.2,"Lubelskie"
"Y15-24","PL32",2002,40,"Podkarpackie"
"Y15-24","PL33",2002,51.3,"Swietokrzyskie"
"Y15-24","PL34",2002,34.4,"Podlaskie"
"Y15-24","PL4",2002,46.3,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2002,40.9,"Wielkopolskie"
"Y15-24","PL42",2002,59.4,"Zachodniopomorskie"
"Y15-24","PL43",2002,45.1,"Lubuskie"
"Y15-24","PL5",2002,46.9,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2002,47.7,"Dolnoslaskie"
"Y15-24","PL52",2002,44.3,"Opolskie"
"Y15-24","PL6",2002,46.6,"Region Pólnocny"
"Y15-24","PL61",2002,45.5,"Kujawsko-Pomorskie"
"Y15-24","PL62",2002,53,"Warminsko-Mazurskie"
"Y15-24","PL63",2002,44.4,"Pomorskie"
"Y15-24","PT",2002,10.5,"Portugal"
"Y15-24","PT1",2002,10.7,"Continente"
"Y15-24","PT11",2002,8.1,"Norte"
"Y15-24","PT15",2002,NA,"Algarve"
"Y15-24","PT16",2002,9.4,"Centro (PT)"
"Y15-24","PT17",2002,15,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2002,NA,"Alentejo"
"Y15-24","PT2",2002,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2002,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2002,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2002,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2002,22.2,"Romania"
"Y15-24","RO1",2002,20.5,"Macroregiunea unu"
"Y15-24","RO11",2002,17.7,"Nord-Vest"
"Y15-24","RO12",2002,23.7,"Centru"
"Y15-24","RO2",2002,20.3,"Macroregiunea doi"
"Y15-24","RO21",2002,17.2,"Nord-Est"
"Y15-24","RO22",2002,25.4,"Sud-Est"
"Y15-24","RO3",2002,28,"Macroregiunea trei"
"Y15-24","RO31",2002,28.8,"Sud - Muntenia"
"Y15-24","RO32",2002,26.4,"Bucuresti - Ilfov"
"Y15-24","RO4",2002,20.7,"Macroregiunea patru"
"Y15-24","RO41",2002,24.2,"Sud-Vest Oltenia"
"Y15-24","RO42",2002,16.1,"Vest"
"Y15-24","SE",2002,12.9,"Sweden"
"Y15-24","SE1",2002,12.2,"Östra Sverige"
"Y15-24","SE11",2002,10.1,"Stockholm"
"Y15-24","SE12",2002,14.7,"Östra Mellansverige"
"Y15-24","SE2",2002,13.5,"Södra Sverige"
"Y15-24","SE21",2002,9.6,"Småland med öarna"
"Y15-24","SE22",2002,16.4,"Sydsverige"
"Y15-24","SE23",2002,13.1,"Västsverige"
"Y15-24","SE3",2002,13.1,"Norra Sverige"
"Y15-24","SE31",2002,13.4,"Norra Mellansverige"
"Y15-24","SE32",2002,15.4,"Mellersta Norrland"
"Y15-24","SE33",2002,11.1,"Övre Norrland"
"Y15-24","SI",2002,14.8,"Slovenia"
"Y15-24","SI0",2002,14.8,"Slovenija"
"Y15-24","SI01",2002,17.4,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2002,11.5,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2002,37.7,"Slovakia"
"Y15-24","SK0",2002,37.7,"Slovensko"
"Y15-24","SK01",2002,20,"Bratislavský kraj"
"Y15-24","SK02",2002,35.1,"Západné Slovensko"
"Y15-24","SK03",2002,39.7,"Stredné Slovensko"
"Y15-24","SK04",2002,45.2,"Východné Slovensko"
"Y15-24","UK",2002,10.9,"United Kingdom"
"Y15-24","UKC",2002,12.1,"North East (UK)"
"Y15-24","UKC1",2002,NA,"Tees Valley and Durham"
"Y15-24","UKC2",2002,12.4,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2002,12.9,"North West (UK)"
"Y15-24","UKD1",2002,NA,"Cumbria"
"Y15-24","UKD3",2002,11.9,"Greater Manchester"
"Y15-24","UKD4",2002,13.6,"Lancashire"
"Y15-24","UKE",2002,12.6,"Yorkshire and The Humber"
"Y15-24","UKE1",2002,19.2,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2002,NA,"North Yorkshire"
"Y15-24","UKE3",2002,10.9,"South Yorkshire"
"Y15-24","UKE4",2002,12.5,"West Yorkshire"
"Y15-24","UKF",2002,8.4,"East Midlands (UK)"
"Y15-24","UKF1",2002,9.9,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2002,NA,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2002,NA,"Lincolnshire"
"Y15-24","UKG",2002,12.5,"West Midlands (UK)"
"Y15-24","UKG1",2002,NA,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2002,9.9,"Shropshire and Staffordshire"
"Y15-24","UKG3",2002,15,"West Midlands"
"Y15-24","UKH",2002,7.5,"East of England"
"Y15-24","UKH1",2002,NA,"East Anglia"
"Y15-24","UKH2",2002,8.7,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2002,9.6,"Essex"
"Y15-24","UKI",2002,12.1,"London"
"Y15-24","UKI1",2002,15.2,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2002,10.1,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2002,8.2,"South East (UK)"
"Y15-24","UKJ1",2002,8.6,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2002,6.2,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2002,8.4,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2002,10.2,"Kent"
"Y15-24","UKK",2002,7.6,"South West (UK)"
"Y15-24","UKK1",2002,6.1,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2002,NA,"Dorset and Somerset"
"Y15-24","UKK3",2002,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2002,NA,"Devon"
"Y15-24","UKL",2002,14.8,"Wales"
"Y15-24","UKL1",2002,13.3,"West Wales and The Valleys"
"Y15-24","UKL2",2002,17.3,"East Wales"
"Y15-24","UKM",2002,13.8,"Scotland"
"Y15-24","UKM2",2002,11.9,"Eastern Scotland"
"Y15-24","UKM3",2002,17.7,"South Western Scotland"
"Y15-24","UKM5",2002,NA,"North Eastern Scotland"
"Y15-24","UKM6",2002,NA,"Highlands and Islands"
"Y15-24","UKN",2002,10.4,"Northern Ireland (UK)"
"Y15-24","UKN0",2002,10.4,"Northern Ireland (UK)"
"Y20-64","AT",2002,4.8,"Austria"
"Y20-64","AT1",2002,6,"Ostösterreich"
"Y20-64","AT11",2002,4.9,"Burgenland (AT)"
"Y20-64","AT12",2002,4.6,"Niederösterreich"
"Y20-64","AT13",2002,7.5,"Wien"
"Y20-64","AT2",2002,5.1,"Südösterreich"
"Y20-64","AT21",2002,4.3,"Kärnten"
"Y20-64","AT22",2002,5.5,"Steiermark"
"Y20-64","AT3",2002,3.1,"Westösterreich"
"Y20-64","AT31",2002,3.7,"Oberösterreich"
"Y20-64","AT32",2002,3.1,"Salzburg"
"Y20-64","AT33",2002,2.3,"Tirol"
"Y20-64","AT34",2002,NA,"Vorarlberg"
"Y20-64","BE",2002,6.8,"Belgium"
"Y20-64","BE1",2002,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2002,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2002,4.6,"Vlaams Gewest"
"Y20-64","BE21",2002,4.8,"Prov. Antwerpen"
"Y20-64","BE22",2002,4.1,"Prov. Limburg (BE)"
"Y20-64","BE23",2002,5.3,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2002,4,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2002,4.3,"Prov. West-Vlaanderen"
"Y20-64","BE3",2002,8.4,"Région wallonne"
"Y20-64","BE31",2002,7.4,"Prov. Brabant Wallon"
"Y20-64","BE32",2002,9.2,"Prov. Hainaut"
"Y20-64","BE33",2002,8.8,"Prov. Liège"
"Y20-64","BE34",2002,NA,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2002,8.1,"Prov. Namur"
"Y20-64","BG",2002,17.6,"Bulgaria"
"Y20-64","BG41",2002,13.2,"Yugozapaden"
"Y20-64","CH",2002,2.8,"Switzerland"
"Y20-64","CH0",2002,2.8,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2002,3.4,"Région lémanique"
"Y20-64","CH02",2002,2.2,"Espace Mittelland"
"Y20-64","CH03",2002,2.5,"Nordwestschweiz"
"Y20-64","CH04",2002,4,"Zürich"
"Y20-64","CH05",2002,2.4,"Ostschweiz"
"Y20-64","CH06",2002,1.7,"Zentralschweiz"
"Y20-64","CH07",2002,3.1,"Ticino"
"Y20-64","CY",2002,3.3,"Cyprus"
"Y20-64","CY0",2002,3.3,"Kypros"
"Y20-64","CY00",2002,3.3,"Kypros"
"Y20-64","CZ",2002,6.7,"Czech Republic"
"Y20-64","CZ0",2002,6.7,"Ceská republika"
"Y20-64","CZ01",2002,3.3,"Praha"
"Y20-64","CZ02",2002,4.6,"Strední Cechy"
"Y20-64","CZ03",2002,4.7,"Jihozápad"
"Y20-64","CZ04",2002,10.3,"Severozápad"
"Y20-64","CZ05",2002,5,"Severovýchod"
"Y20-64","CZ06",2002,6.4,"Jihovýchod"
"Y20-64","CZ07",2002,7.9,"Strední Morava"
"Y20-64","CZ08",2002,12.2,"Moravskoslezsko"
"Y20-64","DE",2002,8.6,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2002,4.4,"Baden-Württemberg"
"Y20-64","DE11",2002,4.3,"Stuttgart"
"Y20-64","DE12",2002,5,"Karlsruhe"
"Y20-64","DE13",2002,4.1,"Freiburg"
"Y20-64","DE14",2002,4.2,"Tübingen"
"Y20-64","DE2",2002,4.6,"Bayern"
"Y20-64","DE21",2002,3.4,"Oberbayern"
"Y20-64","DE22",2002,4.5,"Niederbayern"
"Y20-64","DE23",2002,5.1,"Oberpfalz"
"Y20-64","DE24",2002,7.2,"Oberfranken"
"Y20-64","DE25",2002,5.7,"Mittelfranken"
"Y20-64","DE26",2002,5.4,"Unterfranken"
"Y20-64","DE27",2002,4,"Schwaben"
"Y20-64","DE3",2002,15.7,"Berlin"
"Y20-64","DE30",2002,15.7,"Berlin"
"Y20-64","DE4",2002,17.4,"Brandenburg"
"Y20-64","DE40",2002,17.4,"Brandenburg"
"Y20-64","DE5",2002,9.9,"Bremen"
"Y20-64","DE50",2002,9.9,"Bremen"
"Y20-64","DE6",2002,8.3,"Hamburg"
"Y20-64","DE60",2002,8.3,"Hamburg"
"Y20-64","DE7",2002,5.9,"Hessen"
"Y20-64","DE71",2002,5.5,"Darmstadt"
"Y20-64","DE72",2002,5.4,"Gießen"
"Y20-64","DE73",2002,7.4,"Kassel"
"Y20-64","DE8",2002,20,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2002,20,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2002,7.3,"Niedersachsen"
"Y20-64","DE91",2002,9.1,"Braunschweig"
"Y20-64","DE92",2002,7.4,"Hannover"
"Y20-64","DE93",2002,6.2,"Lüneburg"
"Y20-64","DE94",2002,6.6,"Weser-Ems"
"Y20-64","DEA",2002,7.2,"Nordrhein-Westfalen"
"Y20-64","DEA1",2002,7.4,"Düsseldorf"
"Y20-64","DEA2",2002,6.4,"Köln"
"Y20-64","DEA3",2002,6.8,"Münster"
"Y20-64","DEA4",2002,7.4,"Detmold"
"Y20-64","DEA5",2002,8,"Arnsberg"
"Y20-64","DEB",2002,5.7,"Rheinland-Pfalz"
"Y20-64","DEB1",2002,5.8,"Koblenz"
"Y20-64","DEB2",2002,4.8,"Trier"
"Y20-64","DEB3",2002,5.9,"Rheinhessen-Pfalz"
"Y20-64","DEC",2002,7.7,"Saarland"
"Y20-64","DEC0",2002,7.7,"Saarland"
"Y20-64","DED",2002,18.2,"Sachsen"
"Y20-64","DED2",2002,17.8,"Dresden"
"Y20-64","DEE",2002,19.8,"Sachsen-Anhalt"
"Y20-64","DEE0",2002,19.8,"Sachsen-Anhalt"
"Y20-64","DEF",2002,7.6,"Schleswig-Holstein"
"Y20-64","DEF0",2002,7.6,"Schleswig-Holstein"
"Y20-64","DEG",2002,15.5,"Thüringen"
"Y20-64","DEG0",2002,15.5,"Thüringen"
"Y20-64","DK",2002,4.2,"Denmark"
"Y20-64","DK0",2002,4.2,"Danmark"
"Y20-64","EA17",2002,8.4,"Euro area (17 countries)"
"Y20-64","EA18",2002,8.5,"Euro area (18 countries)"
"Y20-64","EA19",2002,8.5,"Euro area (19 countries)"
"Y20-64","EE",2002,9.7,"Estonia"
"Y20-64","EE0",2002,9.7,"Eesti"
"Y20-64","EE00",2002,9.7,"Eesti"
"Y20-64","EL",2002,9.8,"Greece"
"Y20-64","EL1",2002,10.8,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2002,9.5,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2002,10.8,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2002,13.5,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2002,10.9,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2002,9.4,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2002,11.4,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2002,6.7,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2002,10.7,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2002,9.6,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2002,7.5,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2002,9.2,"Attiki"
"Y20-64","EL30",2002,9.2,"Attiki"
"Y20-64","EL4",2002,9.7,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2002,9.3,"Voreio Aigaio"
"Y20-64","EL42",2002,15.6,"Notio Aigaio"
"Y20-64","EL43",2002,6.7,"Kriti"
"Y20-64","ES",2002,10.7,"Spain"
"Y20-64","ES1",2002,11,"Noroeste (ES)"
"Y20-64","ES11",2002,11.7,"Galicia"
"Y20-64","ES12",2002,10,"Principado de Asturias"
"Y20-64","ES13",2002,9.7,"Cantabria"
"Y20-64","ES2",2002,7.4,"Noreste (ES)"
"Y20-64","ES21",2002,8.9,"País Vasco"
"Y20-64","ES22",2002,4.7,"Comunidad Foral de Navarra"
"Y20-64","ES23",2002,7.6,"La Rioja"
"Y20-64","ES24",2002,5.8,"Aragón"
"Y20-64","ES3",2002,6.8,"Comunidad de Madrid"
"Y20-64","ES30",2002,6.8,"Comunidad de Madrid"
"Y20-64","ES4",2002,11.4,"Centro (ES)"
"Y20-64","ES41",2002,10.4,"Castilla y León"
"Y20-64","ES42",2002,9,"Castilla-la Mancha"
"Y20-64","ES43",2002,18,"Extremadura"
"Y20-64","ES5",2002,9.4,"Este (ES)"
"Y20-64","ES51",2002,9,"Cataluña"
"Y20-64","ES52",2002,10.6,"Comunidad Valenciana"
"Y20-64","ES53",2002,6.4,"Illes Balears"
"Y20-64","ES6",2002,16.8,"Sur (ES)"
"Y20-64","ES61",2002,18.1,"Andalucía"
"Y20-64","ES62",2002,10.3,"Región de Murcia"
"Y20-64","ES63",2002,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2002,NA,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2002,10.6,"Canarias (ES)"
"Y20-64","ES70",2002,10.6,"Canarias (ES)"
"Y20-64","EU15",2002,7.5,"European Union (15 countries)"
"Y20-64","EU27",2002,8.8,"European Union (27 countries)"
"Y20-64","EU28",2002,8.8,"European Union (28 countries)"
"Y20-64","FI",2002,8.4,"Finland"
"Y20-64","FI1",2002,8.5,"Manner-Suomi"
"Y20-64","FI19",2002,8.8,"Länsi-Suomi"
"Y20-64","FI2",2002,NA,"Åland"
"Y20-64","FI20",2002,NA,"Åland"
"Y20-64","FR",2002,8.9,"France"
"Y20-64","FR1",2002,8,"Île de France"
"Y20-64","FR10",2002,8,"Île de France"
"Y20-64","FR2",2002,8.3,"Bassin Parisien"
"Y20-64","FR21",2002,8.7,"Champagne-Ardenne"
"Y20-64","FR22",2002,8.1,"Picardie"
"Y20-64","FR23",2002,9.8,"Haute-Normandie"
"Y20-64","FR24",2002,8.4,"Centre (FR)"
"Y20-64","FR25",2002,7.8,"Basse-Normandie"
"Y20-64","FR26",2002,6.5,"Bourgogne"
"Y20-64","FR3",2002,12.5,"Nord - Pas-de-Calais"
"Y20-64","FR30",2002,12.5,"Nord - Pas-de-Calais"
"Y20-64","FR4",2002,7.3,"Est (FR)"
"Y20-64","FR41",2002,7.6,"Lorraine"
"Y20-64","FR42",2002,6.6,"Alsace"
"Y20-64","FR43",2002,8,"Franche-Comté"
"Y20-64","FR5",2002,7.2,"Ouest (FR)"
"Y20-64","FR51",2002,7.4,"Pays de la Loire"
"Y20-64","FR52",2002,6.7,"Bretagne"
"Y20-64","FR53",2002,7.8,"Poitou-Charentes"
"Y20-64","FR6",2002,8.2,"Sud-Ouest (FR)"
"Y20-64","FR61",2002,9.1,"Aquitaine"
"Y20-64","FR62",2002,7.8,"Midi-Pyrénées"
"Y20-64","FR63",2002,5.9,"Limousin"
"Y20-64","FR7",2002,6.7,"Centre-Est (FR)"
"Y20-64","FR71",2002,6.7,"Rhône-Alpes"
"Y20-64","FR72",2002,6.6,"Auvergne"
"Y20-64","FR8",2002,11.7,"Méditerranée"
"Y20-64","FR81",2002,12.9,"Languedoc-Roussillon"
"Y20-64","FR82",2002,11.1,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2002,NA,"Corse"
"Y20-64","FR9",2002,25.8,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2002,25.4,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2002,22.6,"Martinique (NUTS 2010)"
"Y20-64","FR93",2002,23.7,"Guyane (NUTS 2010)"
"Y20-64","FR94",2002,28.4,"Réunion (NUTS 2010)"
"Y20-64","HR",2002,14.4,"Croatia"
"Y20-64","HR0",2002,14.4,"Hrvatska"
"Y20-64","HU",2002,5.5,"Hungary"
"Y20-64","HU1",2002,3.8,"Közép-Magyarország"
"Y20-64","HU10",2002,3.8,"Közép-Magyarország"
"Y20-64","HU2",2002,5.1,"Dunántúl"
"Y20-64","HU21",2002,4.7,"Közép-Dunántúl"
"Y20-64","HU22",2002,3.5,"Nyugat-Dunántúl"
"Y20-64","HU23",2002,7.6,"Dél-Dunántúl"
"Y20-64","HU3",2002,7.1,"Alföld és Észak"
"Y20-64","HU31",2002,7.9,"Észak-Magyarország"
"Y20-64","HU32",2002,7.6,"Észak-Alföld"
"Y20-64","HU33",2002,5.7,"Dél-Alföld"
"Y20-64","IE",2002,3.9,"Ireland"
"Y20-64","IE0",2002,3.9,"Éire/Ireland"
"Y20-64","IE01",2002,5.1,"Border, Midland and Western"
"Y20-64","IE02",2002,3.6,"Southern and Eastern"
"Y20-64","IS",2002,2.7,"Iceland"
"Y20-64","IS0",2002,2.7,"Ísland"
"Y20-64","IS00",2002,2.7,"Ísland"
"Y20-64","IT",2002,8.8,"Italy"
"Y20-64","ITC",2002,4.3,"Nord-Ovest"
"Y20-64","ITC1",2002,5.4,"Piemonte"
"Y20-64","ITC2",2002,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2002,5.7,"Liguria"
"Y20-64","ITC4",2002,3.5,"Lombardia"
"Y20-64","ITF",2002,17,"Sud"
"Y20-64","ITF1",2002,5.5,"Abruzzo"
"Y20-64","ITF2",2002,12.4,"Molise"
"Y20-64","ITF3",2002,20.2,"Campania"
"Y20-64","ITF4",2002,13,"Puglia"
"Y20-64","ITF5",2002,15.2,"Basilicata"
"Y20-64","ITF6",2002,25,"Calabria"
"Y20-64","ITG",2002,19.4,"Isole"
"Y20-64","ITG1",2002,19.8,"Sicilia"
"Y20-64","ITG2",2002,18.1,"Sardegna"
"Y20-64","ITH",2002,3.5,"Nord-Est"
"Y20-64","ITH1",2002,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2002,3.8,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2002,3.7,"Veneto"
"Y20-64","ITH4",2002,4,"Friuli-Venezia Giulia"
"Y20-64","ITI",2002,6.6,"Centro (IT)"
"Y20-64","ITI1",2002,4.9,"Toscana"
"Y20-64","ITI2",2002,5.3,"Umbria"
"Y20-64","ITI4",2002,8.7,"Lazio"
"Y20-64","LT",2002,13,"Lithuania"
"Y20-64","LT0",2002,13,"Lietuva"
"Y20-64","LT00",2002,13,"Lietuva"
"Y20-64","LU",2002,2.4,"Luxembourg"
"Y20-64","LU0",2002,2.4,"Luxembourg"
"Y20-64","LU00",2002,2.4,"Luxembourg"
"Y20-64","LV",2002,13.5,"Latvia"
"Y20-64","LV0",2002,13.5,"Latvija"
"Y20-64","LV00",2002,13.5,"Latvija"
"Y20-64","MT",2002,5.2,"Malta"
"Y20-64","MT0",2002,5.2,"Malta"
"Y20-64","MT00",2002,5.2,"Malta"
"Y20-64","NL",2002,2.2,"Netherlands"
"Y20-64","NL1",2002,2.3,"Noord-Nederland"
"Y20-64","NL11",2002,2.9,"Groningen"
"Y20-64","NL12",2002,2,"Friesland (NL)"
"Y20-64","NL13",2002,2.1,"Drenthe"
"Y20-64","NL2",2002,2.4,"Oost-Nederland"
"Y20-64","NL21",2002,2.7,"Overijssel"
"Y20-64","NL22",2002,2,"Gelderland"
"Y20-64","NL23",2002,3.6,"Flevoland"
"Y20-64","NL3",2002,2.2,"West-Nederland"
"Y20-64","NL31",2002,1.9,"Utrecht"
"Y20-64","NL32",2002,2.1,"Noord-Holland"
"Y20-64","NL33",2002,2.4,"Zuid-Holland"
"Y20-64","NL34",2002,2,"Zeeland"
"Y20-64","NL4",2002,2.1,"Zuid-Nederland"
"Y20-64","NL41",2002,2.2,"Noord-Brabant"
"Y20-64","NL42",2002,1.9,"Limburg (NL)"
"Y20-64","NO",2002,3.1,"Norway"
"Y20-64","NO0",2002,3.1,"Norge"
"Y20-64","NO01",2002,3.1,"Oslo og Akershus"
"Y20-64","NO02",2002,3,"Hedmark og Oppland"
"Y20-64","NO03",2002,3.3,"Sør-Østlandet"
"Y20-64","NO04",2002,2.6,"Agder og Rogaland"
"Y20-64","NO05",2002,2.5,"Vestlandet"
"Y20-64","NO06",2002,3.8,"Trøndelag"
"Y20-64","NO07",2002,3.4,"Nord-Norge"
"Y20-64","PL",2002,19.7,"Poland"
"Y20-64","PL1",2002,17.9,"Region Centralny"
"Y20-64","PL11",2002,19.8,"Lódzkie"
"Y20-64","PL12",2002,16.7,"Mazowieckie"
"Y20-64","PL2",2002,17.9,"Region Poludniowy"
"Y20-64","PL21",2002,15.4,"Malopolskie"
"Y20-64","PL22",2002,19.7,"Slaskie"
"Y20-64","PL3",2002,17.6,"Region Wschodni"
"Y20-64","PL31",2002,16.7,"Lubelskie"
"Y20-64","PL32",2002,18.6,"Podkarpackie"
"Y20-64","PL33",2002,18.6,"Swietokrzyskie"
"Y20-64","PL34",2002,16.6,"Podlaskie"
"Y20-64","PL4",2002,21.6,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2002,18.4,"Wielkopolskie"
"Y20-64","PL42",2002,25.9,"Zachodniopomorskie"
"Y20-64","PL43",2002,25.5,"Lubuskie"
"Y20-64","PL5",2002,23.7,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2002,24.8,"Dolnoslaskie"
"Y20-64","PL52",2002,20.6,"Opolskie"
"Y20-64","PL6",2002,22.4,"Region Pólnocny"
"Y20-64","PL61",2002,21.9,"Kujawsko-Pomorskie"
"Y20-64","PL62",2002,26.8,"Warminsko-Mazurskie"
"Y20-64","PL63",2002,20.2,"Pomorskie"
"Y20-64","PT",2002,4.5,"Portugal"
"Y20-64","PT1",2002,4.6,"Continente"
"Y20-64","PT11",2002,4.1,"Norte"
"Y20-64","PT15",2002,4.2,"Algarve"
"Y20-64","PT16",2002,2.9,"Centro (PT)"
"Y20-64","PT17",2002,6.1,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2002,6.9,"Alentejo"
"Y20-64","PT2",2002,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2002,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2002,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2002,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2002,8.2,"Romania"
"Y20-64","RO1",2002,7.7,"Macroregiunea unu"
"Y20-64","RO11",2002,7.6,"Nord-Vest"
"Y20-64","RO12",2002,7.8,"Centru"
"Y20-64","RO2",2002,8.5,"Macroregiunea doi"
"Y20-64","RO21",2002,7.3,"Nord-Est"
"Y20-64","RO22",2002,10.2,"Sud-Est"
"Y20-64","RO3",2002,9.5,"Macroregiunea trei"
"Y20-64","RO31",2002,10.4,"Sud - Muntenia"
"Y20-64","RO32",2002,8.3,"Bucuresti - Ilfov"
"Y20-64","RO4",2002,6.5,"Macroregiunea patru"
"Y20-64","RO41",2002,6.7,"Sud-Vest Oltenia"
"Y20-64","RO42",2002,6.2,"Vest"
"Y20-64","SE",2002,4.4,"Sweden"
"Y20-64","SE1",2002,3.9,"Östra Sverige"
"Y20-64","SE11",2002,3.2,"Stockholm"
"Y20-64","SE12",2002,4.8,"Östra Mellansverige"
"Y20-64","SE2",2002,4.3,"Södra Sverige"
"Y20-64","SE21",2002,3.3,"Småland med öarna"
"Y20-64","SE22",2002,5.4,"Sydsverige"
"Y20-64","SE23",2002,4,"Västsverige"
"Y20-64","SE3",2002,5.6,"Norra Sverige"
"Y20-64","SE31",2002,5.6,"Norra Mellansverige"
"Y20-64","SE32",2002,5.6,"Mellersta Norrland"
"Y20-64","SE33",2002,5.7,"Övre Norrland"
"Y20-64","SI",2002,5.9,"Slovenia"
"Y20-64","SI0",2002,5.9,"Slovenija"
"Y20-64","SI01",2002,6.8,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2002,4.8,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2002,17.8,"Slovakia"
"Y20-64","SK0",2002,17.8,"Slovensko"
"Y20-64","SK01",2002,8.3,"Bratislavský kraj"
"Y20-64","SK02",2002,16.6,"Západné Slovensko"
"Y20-64","SK03",2002,20.8,"Stredné Slovensko"
"Y20-64","SK04",2002,21,"Východné Slovensko"
"Y20-64","UK",2002,4.5,"United Kingdom"
"Y20-64","UKC",2002,6,"North East (UK)"
"Y20-64","UKC1",2002,6.1,"Tees Valley and Durham"
"Y20-64","UKC2",2002,6,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2002,4.6,"North West (UK)"
"Y20-64","UKD1",2002,NA,"Cumbria"
"Y20-64","UKD3",2002,4.7,"Greater Manchester"
"Y20-64","UKD4",2002,3.8,"Lancashire"
"Y20-64","UKE",2002,4.5,"Yorkshire and The Humber"
"Y20-64","UKE1",2002,5.6,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2002,3.5,"North Yorkshire"
"Y20-64","UKE3",2002,5,"South Yorkshire"
"Y20-64","UKE4",2002,4.2,"West Yorkshire"
"Y20-64","UKF",2002,3.5,"East Midlands (UK)"
"Y20-64","UKF1",2002,4.1,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2002,2.5,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2002,4.1,"Lincolnshire"
"Y20-64","UKG",2002,4.7,"West Midlands (UK)"
"Y20-64","UKG1",2002,2.6,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2002,3.9,"Shropshire and Staffordshire"
"Y20-64","UKG3",2002,6.3,"West Midlands"
"Y20-64","UKH",2002,3.1,"East of England"
"Y20-64","UKH1",2002,3.2,"East Anglia"
"Y20-64","UKH2",2002,2.6,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2002,3.3,"Essex"
"Y20-64","UKI",2002,6,"London"
"Y20-64","UKI1",2002,8.6,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2002,4.4,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2002,3.4,"South East (UK)"
"Y20-64","UKJ1",2002,3.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2002,3.8,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2002,3.3,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2002,3,"Kent"
"Y20-64","UKK",2002,3.2,"South West (UK)"
"Y20-64","UKK1",2002,2.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2002,3.2,"Dorset and Somerset"
"Y20-64","UKK3",2002,NA,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2002,3.5,"Devon"
"Y20-64","UKL",2002,5.1,"Wales"
"Y20-64","UKL1",2002,4.7,"West Wales and The Valleys"
"Y20-64","UKL2",2002,5.7,"East Wales"
"Y20-64","UKM",2002,5.8,"Scotland"
"Y20-64","UKM2",2002,5.1,"Eastern Scotland"
"Y20-64","UKM3",2002,7.4,"South Western Scotland"
"Y20-64","UKM5",2002,NA,"North Eastern Scotland"
"Y20-64","UKM6",2002,5.1,"Highlands and Islands"
"Y20-64","UKN",2002,5.2,"Northern Ireland (UK)"
"Y20-64","UKN0",2002,5.2,"Northern Ireland (UK)"
"Y_GE15","AT",2002,4.8,"Austria"
"Y_GE15","AT1",2002,6.1,"Ostösterreich"
"Y_GE15","AT11",2002,4.9,"Burgenland (AT)"
"Y_GE15","AT12",2002,4.7,"Niederösterreich"
"Y_GE15","AT13",2002,7.7,"Wien"
"Y_GE15","AT2",2002,5.1,"Südösterreich"
"Y_GE15","AT21",2002,4.4,"Kärnten"
"Y_GE15","AT22",2002,5.5,"Steiermark"
"Y_GE15","AT3",2002,3.2,"Westösterreich"
"Y_GE15","AT31",2002,3.8,"Oberösterreich"
"Y_GE15","AT32",2002,3.2,"Salzburg"
"Y_GE15","AT33",2002,2.4,"Tirol"
"Y_GE15","AT34",2002,2.6,"Vorarlberg"
"Y_GE15","BE",2002,6.9,"Belgium"
"Y_GE15","BE1",2002,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2002,15.8,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2002,4.8,"Vlaams Gewest"
"Y_GE15","BE21",2002,4.8,"Prov. Antwerpen"
"Y_GE15","BE22",2002,4.3,"Prov. Limburg (BE)"
"Y_GE15","BE23",2002,5.6,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2002,4.1,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2002,4.5,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2002,8.5,"Région wallonne"
"Y_GE15","BE31",2002,7.4,"Prov. Brabant Wallon"
"Y_GE15","BE32",2002,9.4,"Prov. Hainaut"
"Y_GE15","BE33",2002,8.7,"Prov. Liège"
"Y_GE15","BE34",2002,5,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2002,8.3,"Prov. Namur"
"Y_GE15","BG",2002,18.1,"Bulgaria"
"Y_GE15","BG41",2002,13.6,"Yugozapaden"
"Y_GE15","CH",2002,2.9,"Switzerland"
"Y_GE15","CH0",2002,2.9,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2002,3.8,"Région lémanique"
"Y_GE15","CH02",2002,2.4,"Espace Mittelland"
"Y_GE15","CH03",2002,2.5,"Nordwestschweiz"
"Y_GE15","CH04",2002,4,"Zürich"
"Y_GE15","CH05",2002,2.4,"Ostschweiz"
"Y_GE15","CH06",2002,1.7,"Zentralschweiz"
"Y_GE15","CH07",2002,3.4,"Ticino"
"Y_GE15","CY",2002,3.3,"Cyprus"
"Y_GE15","CY0",2002,3.3,"Kypros"
"Y_GE15","CY00",2002,3.3,"Kypros"
"Y_GE15","CZ",2002,7,"Czech Republic"
"Y_GE15","CZ0",2002,7,"Ceská republika"
"Y_GE15","CZ01",2002,3.4,"Praha"
"Y_GE15","CZ02",2002,4.8,"Strední Cechy"
"Y_GE15","CZ03",2002,4.8,"Jihozápad"
"Y_GE15","CZ04",2002,11.3,"Severozápad"
"Y_GE15","CZ05",2002,5,"Severovýchod"
"Y_GE15","CZ06",2002,6.7,"Jihovýchod"
"Y_GE15","CZ07",2002,8.5,"Strední Morava"
"Y_GE15","CZ08",2002,12.4,"Moravskoslezsko"
"Y_GE15","DE",2002,8.5,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2002,4.4,"Baden-Württemberg"
"Y_GE15","DE11",2002,4.2,"Stuttgart"
"Y_GE15","DE12",2002,5,"Karlsruhe"
"Y_GE15","DE13",2002,4.2,"Freiburg"
"Y_GE15","DE14",2002,4.1,"Tübingen"
"Y_GE15","DE2",2002,4.5,"Bayern"
"Y_GE15","DE21",2002,3.4,"Oberbayern"
"Y_GE15","DE22",2002,4.4,"Niederbayern"
"Y_GE15","DE23",2002,5,"Oberpfalz"
"Y_GE15","DE24",2002,7,"Oberfranken"
"Y_GE15","DE25",2002,5.6,"Mittelfranken"
"Y_GE15","DE26",2002,5.3,"Unterfranken"
"Y_GE15","DE27",2002,4,"Schwaben"
"Y_GE15","DE3",2002,15.6,"Berlin"
"Y_GE15","DE30",2002,15.6,"Berlin"
"Y_GE15","DE4",2002,16.9,"Brandenburg"
"Y_GE15","DE40",2002,16.9,"Brandenburg"
"Y_GE15","DE5",2002,10,"Bremen"
"Y_GE15","DE50",2002,10,"Bremen"
"Y_GE15","DE6",2002,8.2,"Hamburg"
"Y_GE15","DE60",2002,8.2,"Hamburg"
"Y_GE15","DE7",2002,5.9,"Hessen"
"Y_GE15","DE71",2002,5.5,"Darmstadt"
"Y_GE15","DE72",2002,5.5,"Gießen"
"Y_GE15","DE73",2002,7.4,"Kassel"
"Y_GE15","DE8",2002,19.1,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2002,19.1,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2002,7.2,"Niedersachsen"
"Y_GE15","DE91",2002,9.1,"Braunschweig"
"Y_GE15","DE92",2002,7.3,"Hannover"
"Y_GE15","DE93",2002,6.3,"Lüneburg"
"Y_GE15","DE94",2002,6.4,"Weser-Ems"
"Y_GE15","DEA",2002,7.2,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2002,7.3,"Düsseldorf"
"Y_GE15","DEA2",2002,6.3,"Köln"
"Y_GE15","DEA3",2002,6.8,"Münster"
"Y_GE15","DEA4",2002,7.4,"Detmold"
"Y_GE15","DEA5",2002,8,"Arnsberg"
"Y_GE15","DEB",2002,5.6,"Rheinland-Pfalz"
"Y_GE15","DEB1",2002,5.7,"Koblenz"
"Y_GE15","DEB2",2002,4.6,"Trier"
"Y_GE15","DEB3",2002,5.9,"Rheinhessen-Pfalz"
"Y_GE15","DEC",2002,7.6,"Saarland"
"Y_GE15","DEC0",2002,7.6,"Saarland"
"Y_GE15","DED",2002,17.8,"Sachsen"
"Y_GE15","DED2",2002,17.4,"Dresden"
"Y_GE15","DEE",2002,19.2,"Sachsen-Anhalt"
"Y_GE15","DEE0",2002,19.2,"Sachsen-Anhalt"
"Y_GE15","DEF",2002,7.6,"Schleswig-Holstein"
"Y_GE15","DEF0",2002,7.6,"Schleswig-Holstein"
"Y_GE15","DEG",2002,15.1,"Thüringen"
"Y_GE15","DEG0",2002,15.1,"Thüringen"
"Y_GE15","DK",2002,4.3,"Denmark"
"Y_GE15","DK0",2002,4.3,"Danmark"
"Y_GE15","EA17",2002,8.6,"Euro area (17 countries)"
"Y_GE15","EA18",2002,8.7,"Euro area (18 countries)"
"Y_GE15","EA19",2002,8.7,"Euro area (19 countries)"
"Y_GE15","EE",2002,10,"Estonia"
"Y_GE15","EE0",2002,10,"Eesti"
"Y_GE15","EE00",2002,10,"Eesti"
"Y_GE15","EL",2002,10,"Greece"
"Y_GE15","EL1",2002,10.9,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2002,9.7,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2002,10.9,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2002,13.8,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2002,10.9,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2002,9.5,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2002,11.6,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2002,6.8,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2002,10.8,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2002,9.9,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2002,7.4,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2002,9.4,"Attiki"
"Y_GE15","EL30",2002,9.4,"Attiki"
"Y_GE15","EL4",2002,9.9,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2002,9.8,"Voreio Aigaio"
"Y_GE15","EL42",2002,16,"Notio Aigaio"
"Y_GE15","EL43",2002,6.9,"Kriti"
"Y_GE15","ES",2002,11.1,"Spain"
"Y_GE15","ES1",2002,11.3,"Noroeste (ES)"
"Y_GE15","ES11",2002,12.1,"Galicia"
"Y_GE15","ES12",2002,10.3,"Principado de Asturias"
"Y_GE15","ES13",2002,9.7,"Cantabria"
"Y_GE15","ES2",2002,7.6,"Noreste (ES)"
"Y_GE15","ES21",2002,9.2,"País Vasco"
"Y_GE15","ES22",2002,5.1,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2002,7.8,"La Rioja"
"Y_GE15","ES24",2002,5.9,"Aragón"
"Y_GE15","ES3",2002,7,"Comunidad de Madrid"
"Y_GE15","ES30",2002,7,"Comunidad de Madrid"
"Y_GE15","ES4",2002,11.7,"Centro (ES)"
"Y_GE15","ES41",2002,10.6,"Castilla y León"
"Y_GE15","ES42",2002,9.3,"Castilla-la Mancha"
"Y_GE15","ES43",2002,18.4,"Extremadura"
"Y_GE15","ES5",2002,9.9,"Este (ES)"
"Y_GE15","ES51",2002,9.5,"Cataluña"
"Y_GE15","ES52",2002,11.2,"Comunidad Valenciana"
"Y_GE15","ES53",2002,6.7,"Illes Balears"
"Y_GE15","ES6",2002,17.4,"Sur (ES)"
"Y_GE15","ES61",2002,18.6,"Andalucía"
"Y_GE15","ES62",2002,11.2,"Región de Murcia"
"Y_GE15","ES63",2002,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2002,NA,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2002,11.3,"Canarias (ES)"
"Y_GE15","ES70",2002,11.3,"Canarias (ES)"
"Y_GE15","EU15",2002,7.7,"European Union (15 countries)"
"Y_GE15","EU27",2002,9,"European Union (27 countries)"
"Y_GE15","EU28",2002,9,"European Union (28 countries)"
"Y_GE15","FI",2002,10.4,"Finland"
"Y_GE15","FI1",2002,10.4,"Manner-Suomi"
"Y_GE15","FI19",2002,10.9,"Länsi-Suomi"
"Y_GE15","FI2",2002,NA,"Åland"
"Y_GE15","FI20",2002,NA,"Åland"
"Y_GE15","FR",2002,9.2,"France"
"Y_GE15","FR1",2002,8.1,"Île de France"
"Y_GE15","FR10",2002,8.1,"Île de France"
"Y_GE15","FR2",2002,8.6,"Bassin Parisien"
"Y_GE15","FR21",2002,9.3,"Champagne-Ardenne"
"Y_GE15","FR22",2002,8.5,"Picardie"
"Y_GE15","FR23",2002,10.1,"Haute-Normandie"
"Y_GE15","FR24",2002,8.6,"Centre (FR)"
"Y_GE15","FR25",2002,7.9,"Basse-Normandie"
"Y_GE15","FR26",2002,6.9,"Bourgogne"
"Y_GE15","FR3",2002,13.4,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2002,13.4,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2002,7.5,"Est (FR)"
"Y_GE15","FR41",2002,7.8,"Lorraine"
"Y_GE15","FR42",2002,6.7,"Alsace"
"Y_GE15","FR43",2002,8.3,"Franche-Comté"
"Y_GE15","FR5",2002,7.4,"Ouest (FR)"
"Y_GE15","FR51",2002,7.7,"Pays de la Loire"
"Y_GE15","FR52",2002,6.7,"Bretagne"
"Y_GE15","FR53",2002,8,"Poitou-Charentes"
"Y_GE15","FR6",2002,8.5,"Sud-Ouest (FR)"
"Y_GE15","FR61",2002,9.2,"Aquitaine"
"Y_GE15","FR62",2002,8.1,"Midi-Pyrénées"
"Y_GE15","FR63",2002,6.4,"Limousin"
"Y_GE15","FR7",2002,6.9,"Centre-Est (FR)"
"Y_GE15","FR71",2002,6.9,"Rhône-Alpes"
"Y_GE15","FR72",2002,6.9,"Auvergne"
"Y_GE15","FR8",2002,12,"Méditerranée"
"Y_GE15","FR81",2002,13.1,"Languedoc-Roussillon"
"Y_GE15","FR82",2002,11.4,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2002,NA,"Corse"
"Y_GE15","FR9",2002,26.5,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2002,26,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2002,22.9,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2002,24.4,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2002,29.3,"Réunion (NUTS 2010)"
"Y_GE15","HR",2002,15.1,"Croatia"
"Y_GE15","HR0",2002,15.1,"Hrvatska"
"Y_GE15","HU",2002,5.6,"Hungary"
"Y_GE15","HU1",2002,3.8,"Közép-Magyarország"
"Y_GE15","HU10",2002,3.8,"Közép-Magyarország"
"Y_GE15","HU2",2002,5.3,"Dunántúl"
"Y_GE15","HU21",2002,4.9,"Közép-Dunántúl"
"Y_GE15","HU22",2002,3.7,"Nyugat-Dunántúl"
"Y_GE15","HU23",2002,7.9,"Dél-Dunántúl"
"Y_GE15","HU3",2002,7.3,"Alföld és Észak"
"Y_GE15","HU31",2002,8.2,"Észak-Magyarország"
"Y_GE15","HU32",2002,7.8,"Észak-Alföld"
"Y_GE15","HU33",2002,5.9,"Dél-Alföld"
"Y_GE15","IE",2002,4.2,"Ireland"
"Y_GE15","IE0",2002,4.2,"Éire/Ireland"
"Y_GE15","IE01",2002,5.4,"Border, Midland and Western"
"Y_GE15","IE02",2002,3.8,"Southern and Eastern"
"Y_GE15","IS",2002,3,"Iceland"
"Y_GE15","IS0",2002,3,"Ísland"
"Y_GE15","IS00",2002,3,"Ísland"
"Y_GE15","IT",2002,9.2,"Italy"
"Y_GE15","ITC",2002,4.5,"Nord-Ovest"
"Y_GE15","ITC1",2002,5.5,"Piemonte"
"Y_GE15","ITC2",2002,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2002,6.1,"Liguria"
"Y_GE15","ITC4",2002,3.8,"Lombardia"
"Y_GE15","ITF",2002,17.7,"Sud"
"Y_GE15","ITF1",2002,5.8,"Abruzzo"
"Y_GE15","ITF2",2002,12.6,"Molise"
"Y_GE15","ITF3",2002,21.1,"Campania"
"Y_GE15","ITF4",2002,13.6,"Puglia"
"Y_GE15","ITF5",2002,15.4,"Basilicata"
"Y_GE15","ITF6",2002,25.7,"Calabria"
"Y_GE15","ITG",2002,20.2,"Isole"
"Y_GE15","ITG1",2002,20.7,"Sicilia"
"Y_GE15","ITG2",2002,18.9,"Sardegna"
"Y_GE15","ITH",2002,3.6,"Nord-Est"
"Y_GE15","ITH1",2002,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2002,3.8,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2002,3.8,"Veneto"
"Y_GE15","ITH4",2002,4.1,"Friuli-Venezia Giulia"
"Y_GE15","ITI",2002,6.8,"Centro (IT)"
"Y_GE15","ITI1",2002,5,"Toscana"
"Y_GE15","ITI2",2002,5.5,"Umbria"
"Y_GE15","ITI4",2002,8.9,"Lazio"
"Y_GE15","LT",2002,13,"Lithuania"
"Y_GE15","LT0",2002,13,"Lietuva"
"Y_GE15","LT00",2002,13,"Lietuva"
"Y_GE15","LU",2002,2.6,"Luxembourg"
"Y_GE15","LU0",2002,2.6,"Luxembourg"
"Y_GE15","LU00",2002,2.6,"Luxembourg"
"Y_GE15","LV",2002,13.8,"Latvia"
"Y_GE15","LV0",2002,13.8,"Latvija"
"Y_GE15","LV00",2002,13.8,"Latvija"
"Y_GE15","MT",2002,6.9,"Malta"
"Y_GE15","MT0",2002,6.9,"Malta"
"Y_GE15","MT00",2002,6.9,"Malta"
"Y_GE15","NL",2002,2.6,"Netherlands"
"Y_GE15","NL1",2002,2.9,"Noord-Nederland"
"Y_GE15","NL11",2002,3.5,"Groningen"
"Y_GE15","NL12",2002,2.4,"Friesland (NL)"
"Y_GE15","NL13",2002,2.8,"Drenthe"
"Y_GE15","NL2",2002,2.7,"Oost-Nederland"
"Y_GE15","NL21",2002,2.9,"Overijssel"
"Y_GE15","NL22",2002,2.3,"Gelderland"
"Y_GE15","NL23",2002,4.2,"Flevoland"
"Y_GE15","NL3",2002,2.5,"West-Nederland"
"Y_GE15","NL31",2002,2.3,"Utrecht"
"Y_GE15","NL32",2002,2.4,"Noord-Holland"
"Y_GE15","NL33",2002,2.6,"Zuid-Holland"
"Y_GE15","NL34",2002,2.3,"Zeeland"
"Y_GE15","NL4",2002,2.5,"Zuid-Nederland"
"Y_GE15","NL41",2002,2.5,"Noord-Brabant"
"Y_GE15","NL42",2002,2.4,"Limburg (NL)"
"Y_GE15","NO",2002,4,"Norway"
"Y_GE15","NO0",2002,4,"Norge"
"Y_GE15","NO01",2002,3.9,"Oslo og Akershus"
"Y_GE15","NO02",2002,4.3,"Hedmark og Oppland"
"Y_GE15","NO03",2002,4.2,"Sør-Østlandet"
"Y_GE15","NO04",2002,3.4,"Agder og Rogaland"
"Y_GE15","NO05",2002,3.3,"Vestlandet"
"Y_GE15","NO06",2002,5.1,"Trøndelag"
"Y_GE15","NO07",2002,4.9,"Nord-Norge"
"Y_GE15","PL",2002,19.9,"Poland"
"Y_GE15","PL1",2002,18,"Region Centralny"
"Y_GE15","PL11",2002,20.2,"Lódzkie"
"Y_GE15","PL12",2002,16.7,"Mazowieckie"
"Y_GE15","PL2",2002,18.3,"Region Poludniowy"
"Y_GE15","PL21",2002,15.6,"Malopolskie"
"Y_GE15","PL22",2002,20.3,"Slaskie"
"Y_GE15","PL3",2002,17.3,"Region Wschodni"
"Y_GE15","PL31",2002,16.3,"Lubelskie"
"Y_GE15","PL32",2002,18.2,"Podkarpackie"
"Y_GE15","PL33",2002,18.8,"Swietokrzyskie"
"Y_GE15","PL34",2002,16.1,"Podlaskie"
"Y_GE15","PL4",2002,22.1,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2002,18.7,"Wielkopolskie"
"Y_GE15","PL42",2002,26.7,"Zachodniopomorskie"
"Y_GE15","PL43",2002,25.9,"Lubuskie"
"Y_GE15","PL5",2002,24.1,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2002,25.3,"Dolnoslaskie"
"Y_GE15","PL52",2002,20.9,"Opolskie"
"Y_GE15","PL6",2002,22.9,"Region Pólnocny"
"Y_GE15","PL61",2002,22.3,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2002,27.3,"Warminsko-Mazurskie"
"Y_GE15","PL63",2002,20.9,"Pomorskie"
"Y_GE15","PT",2002,4.5,"Portugal"
"Y_GE15","PT1",2002,4.6,"Continente"
"Y_GE15","PT11",2002,4.1,"Norte"
"Y_GE15","PT15",2002,4.5,"Algarve"
"Y_GE15","PT16",2002,2.8,"Centro (PT)"
"Y_GE15","PT17",2002,6.3,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2002,7.1,"Alentejo"
"Y_GE15","PT2",2002,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2002,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2002,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2002,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2002,8.1,"Romania"
"Y_GE15","RO1",2002,7.9,"Macroregiunea unu"
"Y_GE15","RO11",2002,7.6,"Nord-Vest"
"Y_GE15","RO12",2002,8.2,"Centru"
"Y_GE15","RO2",2002,8.3,"Macroregiunea doi"
"Y_GE15","RO21",2002,6.8,"Nord-Est"
"Y_GE15","RO22",2002,10.4,"Sud-Est"
"Y_GE15","RO3",2002,9.6,"Macroregiunea trei"
"Y_GE15","RO31",2002,10.2,"Sud - Muntenia"
"Y_GE15","RO32",2002,8.6,"Bucuresti - Ilfov"
"Y_GE15","RO4",2002,6.2,"Macroregiunea patru"
"Y_GE15","RO41",2002,6.1,"Sud-Vest Oltenia"
"Y_GE15","RO42",2002,6.3,"Vest"
"Y_GE15","SE",2002,5,"Sweden"
"Y_GE15","SE1",2002,4.4,"Östra Sverige"
"Y_GE15","SE11",2002,3.7,"Stockholm"
"Y_GE15","SE12",2002,5.4,"Östra Mellansverige"
"Y_GE15","SE2",2002,5,"Södra Sverige"
"Y_GE15","SE21",2002,3.8,"Småland med öarna"
"Y_GE15","SE22",2002,6.1,"Sydsverige"
"Y_GE15","SE23",2002,4.8,"Västsverige"
"Y_GE15","SE3",2002,5.9,"Norra Sverige"
"Y_GE15","SE31",2002,5.9,"Norra Mellansverige"
"Y_GE15","SE32",2002,5.8,"Mellersta Norrland"
"Y_GE15","SE33",2002,5.9,"Övre Norrland"
"Y_GE15","SI",2002,5.9,"Slovenia"
"Y_GE15","SI0",2002,5.9,"Slovenija"
"Y_GE15","SI01",2002,6.7,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2002,5,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2002,18.7,"Slovakia"
"Y_GE15","SK0",2002,18.7,"Slovensko"
"Y_GE15","SK01",2002,8.7,"Bratislavský kraj"
"Y_GE15","SK02",2002,17.5,"Západné Slovensko"
"Y_GE15","SK03",2002,21.6,"Stredné Slovensko"
"Y_GE15","SK04",2002,22.3,"Východné Slovensko"
"Y_GE15","UK",2002,5,"United Kingdom"
"Y_GE15","UKC",2002,6.7,"North East (UK)"
"Y_GE15","UKC1",2002,6.5,"Tees Valley and Durham"
"Y_GE15","UKC2",2002,6.9,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2002,5.4,"North West (UK)"
"Y_GE15","UKD1",2002,5.1,"Cumbria"
"Y_GE15","UKD3",2002,5.5,"Greater Manchester"
"Y_GE15","UKD4",2002,4.4,"Lancashire"
"Y_GE15","UKE",2002,5.3,"Yorkshire and The Humber"
"Y_GE15","UKE1",2002,6.9,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2002,4,"North Yorkshire"
"Y_GE15","UKE3",2002,5.2,"South Yorkshire"
"Y_GE15","UKE4",2002,5.1,"West Yorkshire"
"Y_GE15","UKF",2002,4.1,"East Midlands (UK)"
"Y_GE15","UKF1",2002,4.6,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2002,3.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2002,4.5,"Lincolnshire"
"Y_GE15","UKG",2002,5.4,"West Midlands (UK)"
"Y_GE15","UKG1",2002,3.2,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2002,4.4,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2002,7.2,"West Midlands"
"Y_GE15","UKH",2002,3.4,"East of England"
"Y_GE15","UKH1",2002,3.3,"East Anglia"
"Y_GE15","UKH2",2002,3.2,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2002,3.7,"Essex"
"Y_GE15","UKI",2002,6.5,"London"
"Y_GE15","UKI1",2002,8.9,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2002,5,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2002,3.8,"South East (UK)"
"Y_GE15","UKJ1",2002,3.8,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2002,3.9,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2002,3.7,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2002,3.9,"Kent"
"Y_GE15","UKK",2002,3.5,"South West (UK)"
"Y_GE15","UKK1",2002,3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2002,3.4,"Dorset and Somerset"
"Y_GE15","UKK3",2002,4.3,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2002,4.1,"Devon"
"Y_GE15","UKL",2002,5.9,"Wales"
"Y_GE15","UKL1",2002,5.6,"West Wales and The Valleys"
"Y_GE15","UKL2",2002,6.3,"East Wales"
"Y_GE15","UKM",2002,6.7,"Scotland"
"Y_GE15","UKM2",2002,5.7,"Eastern Scotland"
"Y_GE15","UKM3",2002,8.7,"South Western Scotland"
"Y_GE15","UKM5",2002,NA,"North Eastern Scotland"
"Y_GE15","UKM6",2002,5.8,"Highlands and Islands"
"Y_GE15","UKN",2002,5.4,"Northern Ireland (UK)"
"Y_GE15","UKN0",2002,5.4,"Northern Ireland (UK)"
"Y_GE25","AT",2002,4.5,"Austria"
"Y_GE25","AT1",2002,5.7,"Ostösterreich"
"Y_GE25","AT11",2002,4.5,"Burgenland (AT)"
"Y_GE25","AT12",2002,4.4,"Niederösterreich"
"Y_GE25","AT13",2002,7.2,"Wien"
"Y_GE25","AT2",2002,4.7,"Südösterreich"
"Y_GE25","AT21",2002,3.6,"Kärnten"
"Y_GE25","AT22",2002,5.2,"Steiermark"
"Y_GE25","AT3",2002,2.9,"Westösterreich"
"Y_GE25","AT31",2002,3.5,"Oberösterreich"
"Y_GE25","AT32",2002,2.8,"Salzburg"
"Y_GE25","AT33",2002,2.3,"Tirol"
"Y_GE25","AT34",2002,NA,"Vorarlberg"
"Y_GE25","BE",2002,6,"Belgium"
"Y_GE25","BE1",2002,14.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2002,14.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2002,4.1,"Vlaams Gewest"
"Y_GE25","BE21",2002,4.3,"Prov. Antwerpen"
"Y_GE25","BE22",2002,3.7,"Prov. Limburg (BE)"
"Y_GE25","BE23",2002,4.6,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2002,3.3,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2002,4.2,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2002,7.1,"Région wallonne"
"Y_GE25","BE31",2002,5.9,"Prov. Brabant Wallon"
"Y_GE25","BE32",2002,7.4,"Prov. Hainaut"
"Y_GE25","BE33",2002,8,"Prov. Liège"
"Y_GE25","BE34",2002,NA,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2002,7,"Prov. Namur"
"Y_GE25","BG",2002,16.1,"Bulgaria"
"Y_GE25","BG41",2002,12.2,"Yugozapaden"
"Y_GE25","CH",2002,2.5,"Switzerland"
"Y_GE25","CH0",2002,2.5,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2002,3.3,"Région lémanique"
"Y_GE25","CH02",2002,2,"Espace Mittelland"
"Y_GE25","CH03",2002,2.4,"Nordwestschweiz"
"Y_GE25","CH04",2002,3.5,"Zürich"
"Y_GE25","CH05",2002,1.6,"Ostschweiz"
"Y_GE25","CH06",2002,1.5,"Zentralschweiz"
"Y_GE25","CH07",2002,2.9,"Ticino"
"Y_GE25","CY",2002,2.8,"Cyprus"
"Y_GE25","CY0",2002,2.8,"Kypros"
"Y_GE25","CY00",2002,2.8,"Kypros"
"Y_GE25","CZ",2002,6,"Czech Republic"
"Y_GE25","CZ0",2002,6,"Ceská republika"
"Y_GE25","CZ01",2002,2.9,"Praha"
"Y_GE25","CZ02",2002,4.3,"Strední Cechy"
"Y_GE25","CZ03",2002,4.4,"Jihozápad"
"Y_GE25","CZ04",2002,9.2,"Severozápad"
"Y_GE25","CZ05",2002,4.4,"Severovýchod"
"Y_GE25","CZ06",2002,5.6,"Jihovýchod"
"Y_GE25","CZ07",2002,7.1,"Strední Morava"
"Y_GE25","CZ08",2002,10.9,"Moravskoslezsko"
"Y_GE25","DE",2002,8.4,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2002,4.3,"Baden-Württemberg"
"Y_GE25","DE11",2002,4.1,"Stuttgart"
"Y_GE25","DE12",2002,4.8,"Karlsruhe"
"Y_GE25","DE13",2002,4,"Freiburg"
"Y_GE25","DE14",2002,4.1,"Tübingen"
"Y_GE25","DE2",2002,4.5,"Bayern"
"Y_GE25","DE21",2002,3.4,"Oberbayern"
"Y_GE25","DE22",2002,4.2,"Niederbayern"
"Y_GE25","DE23",2002,4.8,"Oberpfalz"
"Y_GE25","DE24",2002,7,"Oberfranken"
"Y_GE25","DE25",2002,5.6,"Mittelfranken"
"Y_GE25","DE26",2002,5.1,"Unterfranken"
"Y_GE25","DE27",2002,3.9,"Schwaben"
"Y_GE25","DE3",2002,15.1,"Berlin"
"Y_GE25","DE30",2002,15.1,"Berlin"
"Y_GE25","DE4",2002,16.9,"Brandenburg"
"Y_GE25","DE40",2002,16.9,"Brandenburg"
"Y_GE25","DE5",2002,9.4,"Bremen"
"Y_GE25","DE50",2002,9.4,"Bremen"
"Y_GE25","DE6",2002,8,"Hamburg"
"Y_GE25","DE60",2002,8,"Hamburg"
"Y_GE25","DE7",2002,5.7,"Hessen"
"Y_GE25","DE71",2002,5.3,"Darmstadt"
"Y_GE25","DE72",2002,5.3,"Gießen"
"Y_GE25","DE73",2002,7.1,"Kassel"
"Y_GE25","DE8",2002,19.9,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2002,19.9,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2002,7,"Niedersachsen"
"Y_GE25","DE91",2002,9,"Braunschweig"
"Y_GE25","DE92",2002,7.1,"Hannover"
"Y_GE25","DE93",2002,5.8,"Lüneburg"
"Y_GE25","DE94",2002,6.3,"Weser-Ems"
"Y_GE25","DEA",2002,7,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2002,7.2,"Düsseldorf"
"Y_GE25","DEA2",2002,6.3,"Köln"
"Y_GE25","DEA3",2002,6.6,"Münster"
"Y_GE25","DEA4",2002,7,"Detmold"
"Y_GE25","DEA5",2002,7.9,"Arnsberg"
"Y_GE25","DEB",2002,5.4,"Rheinland-Pfalz"
"Y_GE25","DEB1",2002,5.4,"Koblenz"
"Y_GE25","DEB2",2002,4.7,"Trier"
"Y_GE25","DEB3",2002,5.5,"Rheinhessen-Pfalz"
"Y_GE25","DEC",2002,7.3,"Saarland"
"Y_GE25","DEC0",2002,7.3,"Saarland"
"Y_GE25","DED",2002,18.2,"Sachsen"
"Y_GE25","DED2",2002,17.5,"Dresden"
"Y_GE25","DEE",2002,19.8,"Sachsen-Anhalt"
"Y_GE25","DEE0",2002,19.8,"Sachsen-Anhalt"
"Y_GE25","DEF",2002,7.3,"Schleswig-Holstein"
"Y_GE25","DEF0",2002,7.3,"Schleswig-Holstein"
"Y_GE25","DEG",2002,15.6,"Thüringen"
"Y_GE25","DEG0",2002,15.6,"Thüringen"
"Y_GE25","DK",2002,3.8,"Denmark"
"Y_GE25","DK0",2002,3.8,"Danmark"
"Y_GE25","EA17",2002,7.6,"Euro area (17 countries)"
"Y_GE25","EA18",2002,7.6,"Euro area (18 countries)"
"Y_GE25","EA19",2002,7.7,"Euro area (19 countries)"
"Y_GE25","EE",2002,8.9,"Estonia"
"Y_GE25","EE0",2002,8.9,"Eesti"
"Y_GE25","EE00",2002,8.9,"Eesti"
"Y_GE25","EL",2002,8,"Greece"
"Y_GE25","EL1",2002,9,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2002,7.7,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2002,9.2,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2002,11.7,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2002,8.6,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2002,7.3,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2002,8.8,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2002,5.6,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2002,8.4,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2002,7.4,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2002,5.8,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2002,7.8,"Attiki"
"Y_GE25","EL30",2002,7.8,"Attiki"
"Y_GE25","EL4",2002,7.4,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2002,7,"Voreio Aigaio"
"Y_GE25","EL42",2002,12.9,"Notio Aigaio"
"Y_GE25","EL43",2002,4.8,"Kriti"
"Y_GE25","ES",2002,9.6,"Spain"
"Y_GE25","ES1",2002,9.8,"Noroeste (ES)"
"Y_GE25","ES11",2002,10.5,"Galicia"
"Y_GE25","ES12",2002,8.9,"Principado de Asturias"
"Y_GE25","ES13",2002,8.3,"Cantabria"
"Y_GE25","ES2",2002,6.6,"Noreste (ES)"
"Y_GE25","ES21",2002,8,"País Vasco"
"Y_GE25","ES22",2002,4.3,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2002,6.9,"La Rioja"
"Y_GE25","ES24",2002,5.1,"Aragón"
"Y_GE25","ES3",2002,6,"Comunidad de Madrid"
"Y_GE25","ES30",2002,6,"Comunidad de Madrid"
"Y_GE25","ES4",2002,10.2,"Centro (ES)"
"Y_GE25","ES41",2002,8.9,"Castilla y León"
"Y_GE25","ES42",2002,8,"Castilla-la Mancha"
"Y_GE25","ES43",2002,17,"Extremadura"
"Y_GE25","ES5",2002,8.3,"Este (ES)"
"Y_GE25","ES51",2002,7.9,"Cataluña"
"Y_GE25","ES52",2002,9.5,"Comunidad Valenciana"
"Y_GE25","ES53",2002,5.6,"Illes Balears"
"Y_GE25","ES6",2002,15.4,"Sur (ES)"
"Y_GE25","ES61",2002,16.6,"Andalucía"
"Y_GE25","ES62",2002,9.2,"Región de Murcia"
"Y_GE25","ES63",2002,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2002,NA,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2002,9.9,"Canarias (ES)"
"Y_GE25","ES70",2002,9.9,"Canarias (ES)"
"Y_GE25","EU15",2002,6.8,"European Union (15 countries)"
"Y_GE25","EU27",2002,7.7,"European Union (27 countries)"
"Y_GE25","EU28",2002,7.8,"European Union (28 countries)"
"Y_GE25","FI",2002,7.3,"Finland"
"Y_GE25","FI1",2002,7.4,"Manner-Suomi"
"Y_GE25","FI19",2002,7.4,"Länsi-Suomi"
"Y_GE25","FI2",2002,NA,"Åland"
"Y_GE25","FI20",2002,NA,"Åland"
"Y_GE25","FR",2002,7.9,"France"
"Y_GE25","FR1",2002,7.5,"Île de France"
"Y_GE25","FR10",2002,7.5,"Île de France"
"Y_GE25","FR2",2002,7.4,"Bassin Parisien"
"Y_GE25","FR21",2002,7.2,"Champagne-Ardenne"
"Y_GE25","FR22",2002,7.1,"Picardie"
"Y_GE25","FR23",2002,8.7,"Haute-Normandie"
"Y_GE25","FR24",2002,7.8,"Centre (FR)"
"Y_GE25","FR25",2002,7,"Basse-Normandie"
"Y_GE25","FR26",2002,5.9,"Bourgogne"
"Y_GE25","FR3",2002,10.8,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2002,10.8,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2002,6.1,"Est (FR)"
"Y_GE25","FR41",2002,6.1,"Lorraine"
"Y_GE25","FR42",2002,5.8,"Alsace"
"Y_GE25","FR43",2002,6.7,"Franche-Comté"
"Y_GE25","FR5",2002,6.3,"Ouest (FR)"
"Y_GE25","FR51",2002,6.7,"Pays de la Loire"
"Y_GE25","FR52",2002,5.7,"Bretagne"
"Y_GE25","FR53",2002,6.9,"Poitou-Charentes"
"Y_GE25","FR6",2002,7.4,"Sud-Ouest (FR)"
"Y_GE25","FR61",2002,8.2,"Aquitaine"
"Y_GE25","FR62",2002,7,"Midi-Pyrénées"
"Y_GE25","FR63",2002,5,"Limousin"
"Y_GE25","FR7",2002,5.8,"Centre-Est (FR)"
"Y_GE25","FR71",2002,5.8,"Rhône-Alpes"
"Y_GE25","FR72",2002,6.2,"Auvergne"
"Y_GE25","FR8",2002,10.6,"Méditerranée"
"Y_GE25","FR81",2002,11.2,"Languedoc-Roussillon"
"Y_GE25","FR82",2002,10.2,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2002,NA,"Corse"
"Y_GE25","FR9",2002,23.4,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2002,23,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2002,20.2,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2002,22,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2002,25.9,"Réunion (NUTS 2010)"
"Y_GE25","HR",2002,12,"Croatia"
"Y_GE25","HR0",2002,12,"Hrvatska"
"Y_GE25","HU",2002,4.9,"Hungary"
"Y_GE25","HU1",2002,3.4,"Közép-Magyarország"
"Y_GE25","HU10",2002,3.4,"Közép-Magyarország"
"Y_GE25","HU2",2002,4.5,"Dunántúl"
"Y_GE25","HU21",2002,4.1,"Közép-Dunántúl"
"Y_GE25","HU22",2002,3.1,"Nyugat-Dunántúl"
"Y_GE25","HU23",2002,6.8,"Dél-Dunántúl"
"Y_GE25","HU3",2002,6.4,"Alföld és Észak"
"Y_GE25","HU31",2002,7,"Észak-Magyarország"
"Y_GE25","HU32",2002,7,"Észak-Alföld"
"Y_GE25","HU33",2002,5.2,"Dél-Alföld"
"Y_GE25","IE",2002,3.5,"Ireland"
"Y_GE25","IE0",2002,3.5,"Éire/Ireland"
"Y_GE25","IE01",2002,4.5,"Border, Midland and Western"
"Y_GE25","IE02",2002,3.1,"Southern and Eastern"
"Y_GE25","IS",2002,2.3,"Iceland"
"Y_GE25","IS0",2002,2.3,"Ísland"
"Y_GE25","IS00",2002,2.3,"Ísland"
"Y_GE25","IT",2002,7.3,"Italy"
"Y_GE25","ITC",2002,3.6,"Nord-Ovest"
"Y_GE25","ITC1",2002,4.5,"Piemonte"
"Y_GE25","ITC2",2002,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2002,4.7,"Liguria"
"Y_GE25","ITC4",2002,3,"Lombardia"
"Y_GE25","ITF",2002,13.9,"Sud"
"Y_GE25","ITF1",2002,4.9,"Abruzzo"
"Y_GE25","ITF2",2002,10.5,"Molise"
"Y_GE25","ITF3",2002,16.1,"Campania"
"Y_GE25","ITF4",2002,10.5,"Puglia"
"Y_GE25","ITF5",2002,12.5,"Basilicata"
"Y_GE25","ITF6",2002,21.5,"Calabria"
"Y_GE25","ITG",2002,16.5,"Isole"
"Y_GE25","ITG1",2002,16.9,"Sicilia"
"Y_GE25","ITG2",2002,15.3,"Sardegna"
"Y_GE25","ITH",2002,3.2,"Nord-Est"
"Y_GE25","ITH1",2002,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2002,3.6,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2002,3.5,"Veneto"
"Y_GE25","ITH4",2002,3.6,"Friuli-Venezia Giulia"
"Y_GE25","ITI",2002,5.4,"Centro (IT)"
"Y_GE25","ITI1",2002,4,"Toscana"
"Y_GE25","ITI2",2002,4.6,"Umbria"
"Y_GE25","ITI4",2002,7,"Lazio"
"Y_GE25","LT",2002,12.2,"Lithuania"
"Y_GE25","LT0",2002,12.2,"Lietuva"
"Y_GE25","LT00",2002,12.2,"Lietuva"
"Y_GE25","LU",2002,2.2,"Luxembourg"
"Y_GE25","LU0",2002,2.2,"Luxembourg"
"Y_GE25","LU00",2002,2.2,"Luxembourg"
"Y_GE25","LV",2002,12.3,"Latvia"
"Y_GE25","LV0",2002,12.3,"Latvija"
"Y_GE25","LV00",2002,12.3,"Latvija"
"Y_GE25","MT",2002,4.5,"Malta"
"Y_GE25","MT0",2002,4.5,"Malta"
"Y_GE25","MT00",2002,4.5,"Malta"
"Y_GE25","NL",2002,2.1,"Netherlands"
"Y_GE25","NL1",2002,2.2,"Noord-Nederland"
"Y_GE25","NL11",2002,2.9,"Groningen"
"Y_GE25","NL12",2002,1.8,"Friesland (NL)"
"Y_GE25","NL13",2002,1.9,"Drenthe"
"Y_GE25","NL2",2002,2.3,"Oost-Nederland"
"Y_GE25","NL21",2002,2.6,"Overijssel"
"Y_GE25","NL22",2002,1.9,"Gelderland"
"Y_GE25","NL23",2002,3.6,"Flevoland"
"Y_GE25","NL3",2002,2.2,"West-Nederland"
"Y_GE25","NL31",2002,1.9,"Utrecht"
"Y_GE25","NL32",2002,2.1,"Noord-Holland"
"Y_GE25","NL33",2002,2.3,"Zuid-Holland"
"Y_GE25","NL34",2002,2.1,"Zeeland"
"Y_GE25","NL4",2002,1.9,"Zuid-Nederland"
"Y_GE25","NL41",2002,2,"Noord-Brabant"
"Y_GE25","NL42",2002,1.8,"Limburg (NL)"
"Y_GE25","NO",2002,2.6,"Norway"
"Y_GE25","NO0",2002,2.6,"Norge"
"Y_GE25","NO01",2002,2.9,"Oslo og Akershus"
"Y_GE25","NO02",2002,2.7,"Hedmark og Oppland"
"Y_GE25","NO03",2002,2.8,"Sør-Østlandet"
"Y_GE25","NO04",2002,1.8,"Agder og Rogaland"
"Y_GE25","NO05",2002,1.8,"Vestlandet"
"Y_GE25","NO06",2002,3.2,"Trøndelag"
"Y_GE25","NO07",2002,3,"Nord-Norge"
"Y_GE25","PL",2002,16.6,"Poland"
"Y_GE25","PL1",2002,15.5,"Region Centralny"
"Y_GE25","PL11",2002,17,"Lódzkie"
"Y_GE25","PL12",2002,14.5,"Mazowieckie"
"Y_GE25","PL2",2002,15,"Region Poludniowy"
"Y_GE25","PL21",2002,12.4,"Malopolskie"
"Y_GE25","PL22",2002,17,"Slaskie"
"Y_GE25","PL3",2002,14.1,"Region Wschodni"
"Y_GE25","PL31",2002,12.9,"Lubelskie"
"Y_GE25","PL32",2002,15.5,"Podkarpackie"
"Y_GE25","PL33",2002,14.2,"Swietokrzyskie"
"Y_GE25","PL34",2002,13.7,"Podlaskie"
"Y_GE25","PL4",2002,18.4,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2002,15.1,"Wielkopolskie"
"Y_GE25","PL42",2002,21.9,"Zachodniopomorskie"
"Y_GE25","PL43",2002,23.2,"Lubuskie"
"Y_GE25","PL5",2002,20.5,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2002,21.6,"Dolnoslaskie"
"Y_GE25","PL52",2002,17.5,"Opolskie"
"Y_GE25","PL6",2002,19.2,"Region Pólnocny"
"Y_GE25","PL61",2002,18.9,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2002,23.7,"Warminsko-Mazurskie"
"Y_GE25","PL63",2002,16.7,"Pomorskie"
"Y_GE25","PT",2002,3.7,"Portugal"
"Y_GE25","PT1",2002,3.8,"Continente"
"Y_GE25","PT11",2002,3.5,"Norte"
"Y_GE25","PT15",2002,NA,"Algarve"
"Y_GE25","PT16",2002,2,"Centro (PT)"
"Y_GE25","PT17",2002,5.2,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2002,6.2,"Alentejo"
"Y_GE25","PT2",2002,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2002,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2002,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2002,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2002,6.1,"Romania"
"Y_GE25","RO1",2002,5.9,"Macroregiunea unu"
"Y_GE25","RO11",2002,5.9,"Nord-Vest"
"Y_GE25","RO12",2002,5.9,"Centru"
"Y_GE25","RO2",2002,6.5,"Macroregiunea doi"
"Y_GE25","RO21",2002,5.2,"Nord-Est"
"Y_GE25","RO22",2002,8.3,"Sud-Est"
"Y_GE25","RO3",2002,7.3,"Macroregiunea trei"
"Y_GE25","RO31",2002,7.7,"Sud - Muntenia"
"Y_GE25","RO32",2002,6.6,"Bucuresti - Ilfov"
"Y_GE25","RO4",2002,4.5,"Macroregiunea patru"
"Y_GE25","RO41",2002,4.1,"Sud-Vest Oltenia"
"Y_GE25","RO42",2002,5.2,"Vest"
"Y_GE25","SE",2002,3.9,"Sweden"
"Y_GE25","SE1",2002,3.5,"Östra Sverige"
"Y_GE25","SE11",2002,3,"Stockholm"
"Y_GE25","SE12",2002,4.1,"Östra Mellansverige"
"Y_GE25","SE2",2002,3.9,"Södra Sverige"
"Y_GE25","SE21",2002,3,"Småland med öarna"
"Y_GE25","SE22",2002,4.7,"Sydsverige"
"Y_GE25","SE23",2002,3.8,"Västsverige"
"Y_GE25","SE3",2002,5,"Norra Sverige"
"Y_GE25","SE31",2002,5.1,"Norra Mellansverige"
"Y_GE25","SE32",2002,4.6,"Mellersta Norrland"
"Y_GE25","SE33",2002,5.2,"Övre Norrland"
"Y_GE25","SI",2002,4.9,"Slovenia"
"Y_GE25","SI0",2002,4.9,"Slovenija"
"Y_GE25","SI01",2002,5.4,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2002,4.3,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2002,15.4,"Slovakia"
"Y_GE25","SK0",2002,15.4,"Slovensko"
"Y_GE25","SK01",2002,7.1,"Bratislavský kraj"
"Y_GE25","SK02",2002,14.4,"Západné Slovensko"
"Y_GE25","SK03",2002,18.3,"Stredné Slovensko"
"Y_GE25","SK04",2002,18.1,"Východné Slovensko"
"Y_GE25","UK",2002,4,"United Kingdom"
"Y_GE25","UKC",2002,5.7,"North East (UK)"
"Y_GE25","UKC1",2002,5.5,"Tees Valley and Durham"
"Y_GE25","UKC2",2002,5.8,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2002,4,"North West (UK)"
"Y_GE25","UKD1",2002,NA,"Cumbria"
"Y_GE25","UKD3",2002,4.2,"Greater Manchester"
"Y_GE25","UKD4",2002,2.8,"Lancashire"
"Y_GE25","UKE",2002,3.9,"Yorkshire and The Humber"
"Y_GE25","UKE1",2002,4.5,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2002,3.5,"North Yorkshire"
"Y_GE25","UKE3",2002,4,"South Yorkshire"
"Y_GE25","UKE4",2002,3.8,"West Yorkshire"
"Y_GE25","UKF",2002,3.4,"East Midlands (UK)"
"Y_GE25","UKF1",2002,3.7,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2002,2.7,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2002,4.2,"Lincolnshire"
"Y_GE25","UKG",2002,4.1,"West Midlands (UK)"
"Y_GE25","UKG1",2002,2.1,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2002,3.4,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2002,5.6,"West Midlands"
"Y_GE25","UKH",2002,2.7,"East of England"
"Y_GE25","UKH1",2002,3.1,"East Anglia"
"Y_GE25","UKH2",2002,2.3,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2002,2.7,"Essex"
"Y_GE25","UKI",2002,5.6,"London"
"Y_GE25","UKI1",2002,7.9,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2002,4.2,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2002,3.1,"South East (UK)"
"Y_GE25","UKJ1",2002,2.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2002,3.6,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2002,2.8,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2002,2.6,"Kent"
"Y_GE25","UKK",2002,2.7,"South West (UK)"
"Y_GE25","UKK1",2002,2.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2002,2.9,"Dorset and Somerset"
"Y_GE25","UKK3",2002,NA,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2002,3.1,"Devon"
"Y_GE25","UKL",2002,4.3,"Wales"
"Y_GE25","UKL1",2002,4.2,"West Wales and The Valleys"
"Y_GE25","UKL2",2002,4.5,"East Wales"
"Y_GE25","UKM",2002,5.3,"Scotland"
"Y_GE25","UKM2",2002,4.7,"Eastern Scotland"
"Y_GE25","UKM3",2002,6.7,"South Western Scotland"
"Y_GE25","UKM5",2002,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2002,4.7,"Highlands and Islands"
"Y_GE25","UKN",2002,4.4,"Northern Ireland (UK)"
"Y_GE25","UKN0",2002,4.4,"Northern Ireland (UK)"
"Y15-24","AT",2001,6,"Austria"
"Y15-24","AT1",2001,6.6,"Ostösterreich"
"Y15-24","AT11",2001,NA,"Burgenland (AT)"
"Y15-24","AT12",2001,5.1,"Niederösterreich"
"Y15-24","AT13",2001,8.5,"Wien"
"Y15-24","AT2",2001,8.7,"Südösterreich"
"Y15-24","AT21",2001,NA,"Kärnten"
"Y15-24","AT22",2001,9.1,"Steiermark"
"Y15-24","AT3",2001,4,"Westösterreich"
"Y15-24","AT31",2001,4.6,"Oberösterreich"
"Y15-24","AT32",2001,NA,"Salzburg"
"Y15-24","AT33",2001,NA,"Tirol"
"Y15-24","AT34",2001,NA,"Vorarlberg"
"Y15-24","BE",2001,15.3,"Belgium"
"Y15-24","BE1",2001,17.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2001,17.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2001,8.7,"Vlaams Gewest"
"Y15-24","BE21",2001,10,"Prov. Antwerpen"
"Y15-24","BE22",2001,13.4,"Prov. Limburg (BE)"
"Y15-24","BE23",2001,8.7,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2001,NA,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2001,NA,"Prov. West-Vlaanderen"
"Y15-24","BE3",2001,27.9,"Région wallonne"
"Y15-24","BE31",2001,NA,"Prov. Brabant Wallon"
"Y15-24","BE32",2001,37.9,"Prov. Hainaut"
"Y15-24","BE33",2001,21.4,"Prov. Liège"
"Y15-24","BE34",2001,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2001,NA,"Prov. Namur"
"Y15-24","BG",2001,39.3,"Bulgaria"
"Y15-24","BG41",2001,31.7,"Yugozapaden"
"Y15-24","CH",2001,5.6,"Switzerland"
"Y15-24","CH0",2001,5.6,"Schweiz/Suisse/Svizzera"
"Y15-24","CH01",2001,13.4,"Région lémanique"
"Y15-24","CH02",2001,4.4,"Espace Mittelland"
"Y15-24","CH03",2001,NA,"Nordwestschweiz"
"Y15-24","CH04",2001,5.9,"Zürich"
"Y15-24","CH05",2001,4.3,"Ostschweiz"
"Y15-24","CH06",2001,NA,"Zentralschweiz"
"Y15-24","CH07",2001,NA,"Ticino"
"Y15-24","CY",2001,8.2,"Cyprus"
"Y15-24","CY0",2001,8.2,"Kypros"
"Y15-24","CY00",2001,8.2,"Kypros"
"Y15-24","CZ",2001,16.3,"Czech Republic"
"Y15-24","CZ0",2001,16.3,"Ceská republika"
"Y15-24","CZ01",2001,9.2,"Praha"
"Y15-24","CZ02",2001,12.7,"Strední Cechy"
"Y15-24","CZ03",2001,7.5,"Jihozápad"
"Y15-24","CZ04",2001,22.1,"Severozápad"
"Y15-24","CZ05",2001,13.2,"Severovýchod"
"Y15-24","CZ06",2001,15.3,"Jihovýchod"
"Y15-24","CZ07",2001,17.9,"Strední Morava"
"Y15-24","CZ08",2001,31.4,"Moravskoslezsko"
"Y15-24","DE",2001,7.8,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2001,3.7,"Baden-Württemberg"
"Y15-24","DE11",2001,4,"Stuttgart"
"Y15-24","DE12",2001,4.1,"Karlsruhe"
"Y15-24","DE13",2001,NA,"Freiburg"
"Y15-24","DE14",2001,NA,"Tübingen"
"Y15-24","DE2",2001,3.8,"Bayern"
"Y15-24","DE21",2001,2.9,"Oberbayern"
"Y15-24","DE22",2001,NA,"Niederbayern"
"Y15-24","DE23",2001,NA,"Oberpfalz"
"Y15-24","DE24",2001,NA,"Oberfranken"
"Y15-24","DE25",2001,5,"Mittelfranken"
"Y15-24","DE26",2001,NA,"Unterfranken"
"Y15-24","DE27",2001,4.4,"Schwaben"
"Y15-24","DE3",2001,17.3,"Berlin"
"Y15-24","DE30",2001,17.3,"Berlin"
"Y15-24","DE4",2001,14.4,"Brandenburg"
"Y15-24","DE40",2001,14.4,"Brandenburg"
"Y15-24","DE5",2001,NA,"Bremen"
"Y15-24","DE50",2001,NA,"Bremen"
"Y15-24","DE6",2001,8.6,"Hamburg"
"Y15-24","DE60",2001,8.6,"Hamburg"
"Y15-24","DE7",2001,5.8,"Hessen"
"Y15-24","DE71",2001,5,"Darmstadt"
"Y15-24","DE72",2001,NA,"Gießen"
"Y15-24","DE73",2001,8.8,"Kassel"
"Y15-24","DE8",2001,13,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2001,13,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2001,7.9,"Niedersachsen"
"Y15-24","DE91",2001,10.5,"Braunschweig"
"Y15-24","DE92",2001,NA,"Hannover"
"Y15-24","DE93",2001,9.8,"Lüneburg"
"Y15-24","DE94",2001,7.6,"Weser-Ems"
"Y15-24","DEA",2001,6.9,"Nordrhein-Westfalen"
"Y15-24","DEA1",2001,6.7,"Düsseldorf"
"Y15-24","DEA2",2001,6.9,"Köln"
"Y15-24","DEA3",2001,6.1,"Münster"
"Y15-24","DEA4",2001,5.2,"Detmold"
"Y15-24","DEA5",2001,8.6,"Arnsberg"
"Y15-24","DEB",2001,6.5,"Rheinland-Pfalz"
"Y15-24","DEC",2001,NA,"Saarland"
"Y15-24","DEC0",2001,NA,"Saarland"
"Y15-24","DED",2001,13.8,"Sachsen"
"Y15-24","DED2",2001,16.5,"Dresden"
"Y15-24","DEE",2001,13.7,"Sachsen-Anhalt"
"Y15-24","DEE0",2001,13.7,"Sachsen-Anhalt"
"Y15-24","DEF",2001,9.4,"Schleswig-Holstein"
"Y15-24","DEF0",2001,9.4,"Schleswig-Holstein"
"Y15-24","DEG",2001,11.7,"Thüringen"
"Y15-24","DEG0",2001,11.7,"Thüringen"
"Y15-24","DK",2001,8.3,"Denmark"
"Y15-24","DK0",2001,8.3,"Danmark"
"Y15-24","EA17",2001,16.1,"Euro area (17 countries)"
"Y15-24","EA18",2001,16.1,"Euro area (18 countries)"
"Y15-24","EA19",2001,16.3,"Euro area (19 countries)"
"Y15-24","EE",2001,24,"Estonia"
"Y15-24","EE0",2001,24,"Eesti"
"Y15-24","EE00",2001,24,"Eesti"
"Y15-24","EL",2001,27.9,"Greece"
"Y15-24","EL1",2001,27.8,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2001,19.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2001,28.3,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2001,38.8,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2001,29.6,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2001,33.5,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2001,36.2,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2001,NA,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2001,33.5,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2001,39.5,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2001,28.9,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2001,27.3,"Attiki"
"Y15-24","EL30",2001,27.3,"Attiki"
"Y15-24","EL4",2001,20.7,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2001,NA,"Voreio Aigaio"
"Y15-24","EL42",2001,20.6,"Notio Aigaio"
"Y15-24","EL43",2001,21,"Kriti"
"Y15-24","ES",2001,20.7,"Spain"
"Y15-24","ES1",2001,22.7,"Noroeste (ES)"
"Y15-24","ES11",2001,25.8,"Galicia"
"Y15-24","ES12",2001,17,"Principado de Asturias"
"Y15-24","ES13",2001,12.6,"Cantabria"
"Y15-24","ES2",2001,15.7,"Noreste (ES)"
"Y15-24","ES21",2001,21.5,"País Vasco"
"Y15-24","ES22",2001,11,"Comunidad Foral de Navarra"
"Y15-24","ES23",2001,NA,"La Rioja"
"Y15-24","ES24",2001,9.2,"Aragón"
"Y15-24","ES3",2001,18,"Comunidad de Madrid"
"Y15-24","ES30",2001,18,"Comunidad de Madrid"
"Y15-24","ES4",2001,21.7,"Centro (ES)"
"Y15-24","ES41",2001,24.1,"Castilla y León"
"Y15-24","ES42",2001,18.9,"Castilla-la Mancha"
"Y15-24","ES43",2001,22.1,"Extremadura"
"Y15-24","ES5",2001,16.4,"Este (ES)"
"Y15-24","ES51",2001,15.8,"Cataluña"
"Y15-24","ES52",2001,17.8,"Comunidad Valenciana"
"Y15-24","ES53",2001,14.5,"Illes Balears"
"Y15-24","ES6",2001,29,"Sur (ES)"
"Y15-24","ES61",2001,31.3,"Andalucía"
"Y15-24","ES62",2001,18.1,"Región de Murcia"
"Y15-24","ES63",2001,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2001,NA,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2001,21.2,"Canarias (ES)"
"Y15-24","ES70",2001,21.2,"Canarias (ES)"
"Y15-24","EU15",2001,14.2,"European Union (15 countries)"
"Y15-24","EU27",2001,17.4,"European Union (27 countries)"
"Y15-24","FI",2001,26.6,"Finland"
"Y15-24","FI1",2001,26.6,"Manner-Suomi"
"Y15-24","FI19",2001,29,"Länsi-Suomi"
"Y15-24","FI2",2001,NA,"Åland"
"Y15-24","FI20",2001,NA,"Åland"
"Y15-24","FR",2001,19,"France"
"Y15-24","FR1",2001,14.1,"Île de France"
"Y15-24","FR10",2001,14.1,"Île de France"
"Y15-24","FR2",2001,18.3,"Bassin Parisien"
"Y15-24","FR21",2001,22.3,"Champagne-Ardenne"
"Y15-24","FR22",2001,23.8,"Picardie"
"Y15-24","FR23",2001,19.8,"Haute-Normandie"
"Y15-24","FR24",2001,16,"Centre (FR)"
"Y15-24","FR25",2001,NA,"Basse-Normandie"
"Y15-24","FR26",2001,NA,"Bourgogne"
"Y15-24","FR3",2001,26.8,"Nord - Pas-de-Calais"
"Y15-24","FR30",2001,26.8,"Nord - Pas-de-Calais"
"Y15-24","FR4",2001,13.6,"Est (FR)"
"Y15-24","FR41",2001,15.3,"Lorraine"
"Y15-24","FR42",2001,13.4,"Alsace"
"Y15-24","FR43",2001,NA,"Franche-Comté"
"Y15-24","FR5",2001,14.1,"Ouest (FR)"
"Y15-24","FR51",2001,15.2,"Pays de la Loire"
"Y15-24","FR52",2001,13,"Bretagne"
"Y15-24","FR53",2001,NA,"Poitou-Charentes"
"Y15-24","FR6",2001,21.4,"Sud-Ouest (FR)"
"Y15-24","FR61",2001,23,"Aquitaine"
"Y15-24","FR62",2001,20.4,"Midi-Pyrénées"
"Y15-24","FR63",2001,NA,"Limousin"
"Y15-24","FR7",2001,15.9,"Centre-Est (FR)"
"Y15-24","FR71",2001,15.2,"Rhône-Alpes"
"Y15-24","FR72",2001,NA,"Auvergne"
"Y15-24","FR8",2001,26.5,"Méditerranée"
"Y15-24","FR81",2001,30.8,"Languedoc-Roussillon"
"Y15-24","FR82",2001,24.1,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2001,NA,"Corse"
"Y15-24","FR9",2001,53.6,"Départements d'outre-mer (NUTS 2010)"
"Y15-24","FR91",2001,56.2,"Guadeloupe (NUTS 2010)"
"Y15-24","FR92",2001,50.3,"Martinique (NUTS 2010)"
"Y15-24","FR93",2001,50.8,"Guyane (NUTS 2010)"
"Y15-24","FR94",2001,54.3,"Réunion (NUTS 2010)"
"Y15-24","HU",2001,10.7,"Hungary"
"Y15-24","HU1",2001,8.8,"Közép-Magyarország"
"Y15-24","HU10",2001,8.8,"Közép-Magyarország"
"Y15-24","HU2",2001,9.7,"Dunántúl"
"Y15-24","HU21",2001,5.3,"Közép-Dunántúl"
"Y15-24","HU22",2001,9.6,"Nyugat-Dunántúl"
"Y15-24","HU23",2001,15.2,"Dél-Dunántúl"
"Y15-24","HU3",2001,12.8,"Alföld és Észak"
"Y15-24","HU31",2001,13.5,"Észak-Magyarország"
"Y15-24","HU32",2001,13.1,"Észak-Alföld"
"Y15-24","HU33",2001,11.8,"Dél-Alföld"
"Y15-24","IE",2001,6.2,"Ireland"
"Y15-24","IE0",2001,6.2,"Éire/Ireland"
"Y15-24","IE01",2001,7.7,"Border, Midland and Western"
"Y15-24","IE02",2001,5.7,"Southern and Eastern"
"Y15-24","IS",2001,5.1,"Iceland"
"Y15-24","IS0",2001,5.1,"Ísland"
"Y15-24","IS00",2001,5.1,"Ísland"
"Y15-24","IT",2001,27.8,"Italy"
"Y15-24","ITC",2001,13.1,"Nord-Ovest"
"Y15-24","ITC1",2001,14.7,"Piemonte"
"Y15-24","ITC2",2001,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2001,25.4,"Liguria"
"Y15-24","ITC4",2001,11.2,"Lombardia"
"Y15-24","ITF",2001,49.2,"Sud"
"Y15-24","ITF1",2001,18.6,"Abruzzo"
"Y15-24","ITF2",2001,38,"Molise"
"Y15-24","ITF3",2001,60.2,"Campania"
"Y15-24","ITF4",2001,37.7,"Puglia"
"Y15-24","ITF5",2001,42.7,"Basilicata"
"Y15-24","ITF6",2001,58.8,"Calabria"
"Y15-24","ITG",2001,51.9,"Isole"
"Y15-24","ITG1",2001,51.8,"Sicilia"
"Y15-24","ITG2",2001,52.1,"Sardegna"
"Y15-24","ITH",2001,8.6,"Nord-Est"
"Y15-24","ITH1",2001,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2001,NA,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2001,7.2,"Veneto"
"Y15-24","ITH4",2001,NA,"Friuli-Venezia Giulia"
"Y15-24","ITI",2001,23.5,"Centro (IT)"
"Y15-24","ITI1",2001,17.3,"Toscana"
"Y15-24","ITI2",2001,NA,"Umbria"
"Y15-24","ITI4",2001,33.4,"Lazio"
"Y15-24","LT",2001,31.6,"Lithuania"
"Y15-24","LT0",2001,31.6,"Lietuva"
"Y15-24","LT00",2001,31.6,"Lietuva"
"Y15-24","LU",2001,6.3,"Luxembourg"
"Y15-24","LU0",2001,6.3,"Luxembourg"
"Y15-24","LU00",2001,6.3,"Luxembourg"
"Y15-24","LV",2001,24.2,"Latvia"
"Y15-24","LV0",2001,24.2,"Latvija"
"Y15-24","LV00",2001,24.2,"Latvija"
"Y15-24","MT",2001,17.6,"Malta"
"Y15-24","MT0",2001,17.6,"Malta"
"Y15-24","MT00",2001,17.6,"Malta"
"Y15-24","NL",2001,4.4,"Netherlands"
"Y15-24","NL1",2001,7,"Noord-Nederland"
"Y15-24","NL11",2001,7.3,"Groningen"
"Y15-24","NL12",2001,7.3,"Friesland (NL)"
"Y15-24","NL13",2001,6.3,"Drenthe"
"Y15-24","NL2",2001,4.1,"Oost-Nederland"
"Y15-24","NL21",2001,5.6,"Overijssel"
"Y15-24","NL22",2001,3.4,"Gelderland"
"Y15-24","NL23",2001,NA,"Flevoland"
"Y15-24","NL3",2001,3.9,"West-Nederland"
"Y15-24","NL31",2001,2,"Utrecht"
"Y15-24","NL32",2001,5,"Noord-Holland"
"Y15-24","NL33",2001,4,"Zuid-Holland"
"Y15-24","NL34",2001,NA,"Zeeland"
"Y15-24","NL4",2001,4.4,"Zuid-Nederland"
"Y15-24","NL41",2001,4,"Noord-Brabant"
"Y15-24","NL42",2001,5.3,"Limburg (NL)"
"Y15-24","NO",2001,12.2,"Norway"
"Y15-24","NO0",2001,12.2,"Norge"
"Y15-24","NO01",2001,6.9,"Oslo og Akershus"
"Y15-24","NO02",2001,13.1,"Hedmark og Oppland"
"Y15-24","NO03",2001,12,"Sør-Østlandet"
"Y15-24","NO04",2001,13.2,"Agder og Rogaland"
"Y15-24","NO05",2001,11.7,"Vestlandet"
"Y15-24","NO06",2001,12.8,"Trøndelag"
"Y15-24","NO07",2001,21.7,"Nord-Norge"
"Y15-24","PL",2001,39.2,"Poland"
"Y15-24","PL1",2001,35.3,"Region Centralny"
"Y15-24","PL11",2001,41.1,"Lódzkie"
"Y15-24","PL12",2001,31.5,"Mazowieckie"
"Y15-24","PL2",2001,37.4,"Region Poludniowy"
"Y15-24","PL21",2001,33.6,"Malopolskie"
"Y15-24","PL22",2001,40.6,"Slaskie"
"Y15-24","PL3",2001,41.3,"Region Wschodni"
"Y15-24","PL31",2001,36.1,"Lubelskie"
"Y15-24","PL32",2001,44.7,"Podkarpackie"
"Y15-24","PL33",2001,49.1,"Swietokrzyskie"
"Y15-24","PL34",2001,37.7,"Podlaskie"
"Y15-24","PL4",2001,41.3,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2001,38.5,"Wielkopolskie"
"Y15-24","PL42",2001,44.6,"Zachodniopomorskie"
"Y15-24","PL43",2001,47.4,"Lubuskie"
"Y15-24","PL5",2001,43.7,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2001,44,"Dolnoslaskie"
"Y15-24","PL52",2001,43,"Opolskie"
"Y15-24","PL6",2001,39.1,"Region Pólnocny"
"Y15-24","PL61",2001,40.1,"Kujawsko-Pomorskie"
"Y15-24","PL62",2001,47.9,"Warminsko-Mazurskie"
"Y15-24","PL63",2001,32.6,"Pomorskie"
"Y15-24","PT",2001,8.9,"Portugal"
"Y15-24","PT1",2001,9.1,"Continente"
"Y15-24","PT11",2001,6.2,"Norte"
"Y15-24","PT15",2001,NA,"Algarve"
"Y15-24","PT16",2001,9.5,"Centro (PT)"
"Y15-24","PT17",2001,12.6,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2001,NA,"Alentejo"
"Y15-24","PT2",2001,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2001,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2001,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2001,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2001,17.6,"Romania"
"Y15-24","RO1",2001,14.9,"Macroregiunea unu"
"Y15-24","RO11",2001,13,"Nord-Vest"
"Y15-24","RO12",2001,17.2,"Centru"
"Y15-24","RO2",2001,18,"Macroregiunea doi"
"Y15-24","RO21",2001,15,"Nord-Est"
"Y15-24","RO22",2001,23.1,"Sud-Est"
"Y15-24","RO3",2001,23.2,"Macroregiunea trei"
"Y15-24","RO31",2001,22.9,"Sud - Muntenia"
"Y15-24","RO32",2001,23.9,"Bucuresti - Ilfov"
"Y15-24","RO4",2001,14.3,"Macroregiunea patru"
"Y15-24","RO41",2001,16.8,"Sud-Vest Oltenia"
"Y15-24","RO42",2001,10.9,"Vest"
"Y15-24","SE",2001,11.7,"Sweden"
"Y15-24","SE1",2001,10.9,"Östra Sverige"
"Y15-24","SE11",2001,8.7,"Stockholm"
"Y15-24","SE12",2001,13.8,"Östra Mellansverige"
"Y15-24","SE2",2001,11.5,"Södra Sverige"
"Y15-24","SE21",2001,7.9,"Småland med öarna"
"Y15-24","SE22",2001,14.7,"Sydsverige"
"Y15-24","SE23",2001,11,"Västsverige"
"Y15-24","SE3",2001,13.8,"Norra Sverige"
"Y15-24","SE31",2001,16.2,"Norra Mellansverige"
"Y15-24","SE32",2001,NA,"Mellersta Norrland"
"Y15-24","SE33",2001,12,"Övre Norrland"
"Y15-24","SI",2001,15.7,"Slovenia"
"Y15-24","SI0",2001,15.7,"Slovenija"
"Y15-24","SI01",2001,17.7,"Vzhodna Slovenija (NUTS 2010)"
"Y15-24","SI02",2001,13.3,"Zahodna Slovenija (NUTS 2010)"
"Y15-24","SK",2001,38.9,"Slovakia"
"Y15-24","SK0",2001,38.9,"Slovensko"
"Y15-24","SK01",2001,19.9,"Bratislavský kraj"
"Y15-24","SK02",2001,35.6,"Západné Slovensko"
"Y15-24","SK03",2001,41.2,"Stredné Slovensko"
"Y15-24","SK04",2001,48.3,"Východné Slovensko"
"Y15-24","UK",2001,10.3,"United Kingdom"
"Y15-24","UKC",2001,13.5,"North East (UK)"
"Y15-24","UKC1",2001,NA,"Tees Valley and Durham"
"Y15-24","UKC2",2001,14.8,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2001,12.9,"North West (UK)"
"Y15-24","UKD1",2001,NA,"Cumbria"
"Y15-24","UKD3",2001,10.8,"Greater Manchester"
"Y15-24","UKD4",2001,NA,"Lancashire"
"Y15-24","UKE",2001,9.8,"Yorkshire and The Humber"
"Y15-24","UKE1",2001,NA,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2001,NA,"North Yorkshire"
"Y15-24","UKE3",2001,NA,"South Yorkshire"
"Y15-24","UKE4",2001,10.3,"West Yorkshire"
"Y15-24","UKF",2001,10.8,"East Midlands (UK)"
"Y15-24","UKF1",2001,13.2,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2001,NA,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2001,NA,"Lincolnshire"
"Y15-24","UKG",2001,9.4,"West Midlands (UK)"
"Y15-24","UKG1",2001,NA,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2001,NA,"Shropshire and Staffordshire"
"Y15-24","UKG3",2001,12.6,"West Midlands"
"Y15-24","UKH",2001,8.5,"East of England"
"Y15-24","UKH1",2001,10.3,"East Anglia"
"Y15-24","UKH2",2001,NA,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2001,NA,"Essex"
"Y15-24","UKI",2001,12.3,"London"
"Y15-24","UKI1",2001,15.5,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2001,10.2,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2001,6.6,"South East (UK)"
"Y15-24","UKJ1",2001,6.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2001,6.4,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2001,NA,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2001,NA,"Kent"
"Y15-24","UKK",2001,6.6,"South West (UK)"
"Y15-24","UKK1",2001,NA,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2001,NA,"Dorset and Somerset"
"Y15-24","UKK3",2001,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2001,NA,"Devon"
"Y15-24","UKL",2001,13.6,"Wales"
"Y15-24","UKL1",2001,15.4,"West Wales and The Valleys"
"Y15-24","UKL2",2001,NA,"East Wales"
"Y15-24","UKM",2001,13.3,"Scotland"
"Y15-24","UKM2",2001,12,"Eastern Scotland"
"Y15-24","UKM3",2001,13.2,"South Western Scotland"
"Y15-24","UKM5",2001,NA,"North Eastern Scotland"
"Y15-24","UKM6",2001,NA,"Highlands and Islands"
"Y15-24","UKN",2001,9.7,"Northern Ireland (UK)"
"Y15-24","UKN0",2001,9.7,"Northern Ireland (UK)"
"Y20-64","AT",2001,3.9,"Austria"
"Y20-64","AT1",2001,4.6,"Ostösterreich"
"Y20-64","AT11",2001,4.9,"Burgenland (AT)"
"Y20-64","AT12",2001,3.2,"Niederösterreich"
"Y20-64","AT13",2001,5.9,"Wien"
"Y20-64","AT2",2001,4.3,"Südösterreich"
"Y20-64","AT21",2001,4.7,"Kärnten"
"Y20-64","AT22",2001,4.1,"Steiermark"
"Y20-64","AT3",2001,2.8,"Westösterreich"
"Y20-64","AT31",2001,3,"Oberösterreich"
"Y20-64","AT32",2001,2,"Salzburg"
"Y20-64","AT33",2001,2.8,"Tirol"
"Y20-64","AT34",2001,2.9,"Vorarlberg"
"Y20-64","BE",2001,6,"Belgium"
"Y20-64","BE1",2001,13,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2001,13,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2001,3.4,"Vlaams Gewest"
"Y20-64","BE21",2001,4.4,"Prov. Antwerpen"
"Y20-64","BE22",2001,3.2,"Prov. Limburg (BE)"
"Y20-64","BE23",2001,3.4,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2001,3.5,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2001,2,"Prov. West-Vlaanderen"
"Y20-64","BE3",2001,9,"Région wallonne"
"Y20-64","BE31",2001,5.6,"Prov. Brabant Wallon"
"Y20-64","BE32",2001,11.3,"Prov. Hainaut"
"Y20-64","BE33",2001,9.2,"Prov. Liège"
"Y20-64","BE34",2001,5.5,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2001,7.5,"Prov. Namur"
"Y20-64","BG",2001,19.3,"Bulgaria"
"Y20-64","BG41",2001,14.9,"Yugozapaden"
"Y20-64","CH",2001,2.2,"Switzerland"
"Y20-64","CH0",2001,2.2,"Schweiz/Suisse/Svizzera"
"Y20-64","CH01",2001,3.1,"Région lémanique"
"Y20-64","CH02",2001,1.6,"Espace Mittelland"
"Y20-64","CH03",2001,2.3,"Nordwestschweiz"
"Y20-64","CH04",2001,2.2,"Zürich"
"Y20-64","CH05",2001,1.6,"Ostschweiz"
"Y20-64","CH06",2001,2.1,"Zentralschweiz"
"Y20-64","CH07",2001,2.8,"Ticino"
"Y20-64","CY",2001,3.8,"Cyprus"
"Y20-64","CY0",2001,3.8,"Kypros"
"Y20-64","CY00",2001,3.8,"Kypros"
"Y20-64","CZ",2001,7.6,"Czech Republic"
"Y20-64","CZ0",2001,7.6,"Ceská republika"
"Y20-64","CZ01",2001,3.7,"Praha"
"Y20-64","CZ02",2001,6.4,"Strední Cechy"
"Y20-64","CZ03",2001,4.9,"Jihozápad"
"Y20-64","CZ04",2001,11.2,"Severozápad"
"Y20-64","CZ05",2001,5.5,"Severovýchod"
"Y20-64","CZ06",2001,6.9,"Jihovýchod"
"Y20-64","CZ07",2001,9,"Strední Morava"
"Y20-64","CZ08",2001,14.3,"Moravskoslezsko"
"Y20-64","DE",2001,7.9,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2001,3.9,"Baden-Württemberg"
"Y20-64","DE11",2001,3.6,"Stuttgart"
"Y20-64","DE12",2001,4.3,"Karlsruhe"
"Y20-64","DE13",2001,4,"Freiburg"
"Y20-64","DE14",2001,3.5,"Tübingen"
"Y20-64","DE2",2001,3.9,"Bayern"
"Y20-64","DE21",2001,2.8,"Oberbayern"
"Y20-64","DE22",2001,3.8,"Niederbayern"
"Y20-64","DE23",2001,4.8,"Oberpfalz"
"Y20-64","DE24",2001,5.5,"Oberfranken"
"Y20-64","DE25",2001,4.9,"Mittelfranken"
"Y20-64","DE26",2001,4.4,"Unterfranken"
"Y20-64","DE27",2001,3.8,"Schwaben"
"Y20-64","DE3",2001,15,"Berlin"
"Y20-64","DE30",2001,15,"Berlin"
"Y20-64","DE4",2001,17.4,"Brandenburg"
"Y20-64","DE40",2001,17.4,"Brandenburg"
"Y20-64","DE5",2001,8.6,"Bremen"
"Y20-64","DE50",2001,8.6,"Bremen"
"Y20-64","DE6",2001,7,"Hamburg"
"Y20-64","DE60",2001,7,"Hamburg"
"Y20-64","DE7",2001,5.5,"Hessen"
"Y20-64","DE71",2001,5.2,"Darmstadt"
"Y20-64","DE72",2001,5.2,"Gießen"
"Y20-64","DE73",2001,6.9,"Kassel"
"Y20-64","DE8",2001,19.3,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2001,19.3,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2001,6.3,"Niedersachsen"
"Y20-64","DE91",2001,8.1,"Braunschweig"
"Y20-64","DE92",2001,6.6,"Hannover"
"Y20-64","DE93",2001,5.8,"Lüneburg"
"Y20-64","DE94",2001,5.3,"Weser-Ems"
"Y20-64","DEA",2001,6.1,"Nordrhein-Westfalen"
"Y20-64","DEA1",2001,6.1,"Düsseldorf"
"Y20-64","DEA2",2001,5.7,"Köln"
"Y20-64","DEA3",2001,5.7,"Münster"
"Y20-64","DEA4",2001,5.9,"Detmold"
"Y20-64","DEA5",2001,6.9,"Arnsberg"
"Y20-64","DEB",2001,5,"Rheinland-Pfalz"
"Y20-64","DEC",2001,5.9,"Saarland"
"Y20-64","DEC0",2001,5.9,"Saarland"
"Y20-64","DED",2001,17.6,"Sachsen"
"Y20-64","DED2",2001,17.8,"Dresden"
"Y20-64","DEE",2001,20.5,"Sachsen-Anhalt"
"Y20-64","DEE0",2001,20.5,"Sachsen-Anhalt"
"Y20-64","DEF",2001,6.4,"Schleswig-Holstein"
"Y20-64","DEF0",2001,6.4,"Schleswig-Holstein"
"Y20-64","DEG",2001,14.3,"Thüringen"
"Y20-64","DEG0",2001,14.3,"Thüringen"
"Y20-64","DK",2001,4,"Denmark"
"Y20-64","DK0",2001,4,"Danmark"
"Y20-64","EA17",2001,8.1,"Euro area (17 countries)"
"Y20-64","EA18",2001,8.1,"Euro area (18 countries)"
"Y20-64","EA19",2001,8.2,"Euro area (19 countries)"
"Y20-64","EE",2001,12.6,"Estonia"
"Y20-64","EE0",2001,12.6,"Eesti"
"Y20-64","EE00",2001,12.6,"Eesti"
"Y20-64","EL",2001,10.2,"Greece"
"Y20-64","EL1",2001,11.1,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2001,9,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2001,10.6,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2001,15.9,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2001,12.2,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2001,10.5,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2001,12.7,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2001,7.6,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2001,9.8,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2001,13.3,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2001,8.6,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2001,10,"Attiki"
"Y20-64","EL30",2001,10,"Attiki"
"Y20-64","EL4",2001,7.2,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2001,6.4,"Voreio Aigaio"
"Y20-64","EL42",2001,9.6,"Notio Aigaio"
"Y20-64","EL43",2001,6.3,"Kriti"
"Y20-64","ES",2001,9.8,"Spain"
"Y20-64","ES1",2001,10,"Noroeste (ES)"
"Y20-64","ES11",2001,11.1,"Galicia"
"Y20-64","ES12",2001,7.8,"Principado de Asturias"
"Y20-64","ES13",2001,8,"Cantabria"
"Y20-64","ES2",2001,7,"Noreste (ES)"
"Y20-64","ES21",2001,9.2,"País Vasco"
"Y20-64","ES22",2001,4.1,"Comunidad Foral de Navarra"
"Y20-64","ES23",2001,4.1,"La Rioja"
"Y20-64","ES24",2001,4.9,"Aragón"
"Y20-64","ES3",2001,6.9,"Comunidad de Madrid"
"Y20-64","ES30",2001,6.9,"Comunidad de Madrid"
"Y20-64","ES4",2001,10,"Centro (ES)"
"Y20-64","ES41",2001,9.3,"Castilla y León"
"Y20-64","ES42",2001,8.9,"Castilla-la Mancha"
"Y20-64","ES43",2001,13.5,"Extremadura"
"Y20-64","ES5",2001,8,"Este (ES)"
"Y20-64","ES51",2001,7.8,"Cataluña"
"Y20-64","ES52",2001,9,"Comunidad Valenciana"
"Y20-64","ES53",2001,5.3,"Illes Balears"
"Y20-64","ES6",2001,16.1,"Sur (ES)"
"Y20-64","ES61",2001,17.6,"Andalucía"
"Y20-64","ES62",2001,8.6,"Región de Murcia"
"Y20-64","ES63",2001,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2001,NA,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2001,9.9,"Canarias (ES)"
"Y20-64","ES70",2001,9.9,"Canarias (ES)"
"Y20-64","EU15",2001,7.1,"European Union (15 countries)"
"Y20-64","EU27",2001,8.4,"European Union (27 countries)"
"Y20-64","FI",2001,8.6,"Finland"
"Y20-64","FI1",2001,8.6,"Manner-Suomi"
"Y20-64","FI19",2001,9.3,"Länsi-Suomi"
"Y20-64","FI2",2001,NA,"Åland"
"Y20-64","FI20",2001,NA,"Åland"
"Y20-64","FR",2001,8.8,"France"
"Y20-64","FR1",2001,7.2,"Île de France"
"Y20-64","FR10",2001,7.2,"Île de France"
"Y20-64","FR2",2001,7.9,"Bassin Parisien"
"Y20-64","FR21",2001,9.6,"Champagne-Ardenne"
"Y20-64","FR22",2001,8.9,"Picardie"
"Y20-64","FR23",2001,8.4,"Haute-Normandie"
"Y20-64","FR24",2001,7,"Centre (FR)"
"Y20-64","FR25",2001,7,"Basse-Normandie"
"Y20-64","FR26",2001,6.9,"Bourgogne"
"Y20-64","FR3",2001,13.2,"Nord - Pas-de-Calais"
"Y20-64","FR30",2001,13.2,"Nord - Pas-de-Calais"
"Y20-64","FR4",2001,6.2,"Est (FR)"
"Y20-64","FR41",2001,7.3,"Lorraine"
"Y20-64","FR42",2001,5.8,"Alsace"
"Y20-64","FR43",2001,4.7,"Franche-Comté"
"Y20-64","FR5",2001,7.2,"Ouest (FR)"
"Y20-64","FR51",2001,7.6,"Pays de la Loire"
"Y20-64","FR52",2001,6.2,"Bretagne"
"Y20-64","FR53",2001,8.5,"Poitou-Charentes"
"Y20-64","FR6",2001,9.1,"Sud-Ouest (FR)"
"Y20-64","FR61",2001,10,"Aquitaine"
"Y20-64","FR62",2001,8.6,"Midi-Pyrénées"
"Y20-64","FR63",2001,7,"Limousin"
"Y20-64","FR7",2001,7,"Centre-Est (FR)"
"Y20-64","FR71",2001,7,"Rhône-Alpes"
"Y20-64","FR72",2001,7.3,"Auvergne"
"Y20-64","FR8",2001,12.5,"Méditerranée"
"Y20-64","FR81",2001,13,"Languedoc-Roussillon"
"Y20-64","FR82",2001,12.2,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2001,NA,"Corse"
"Y20-64","FR9",2001,27,"Départements d'outre-mer (NUTS 2010)"
"Y20-64","FR91",2001,24.8,"Guadeloupe (NUTS 2010)"
"Y20-64","FR92",2001,23.6,"Martinique (NUTS 2010)"
"Y20-64","FR93",2001,27.4,"Guyane (NUTS 2010)"
"Y20-64","FR94",2001,30.2,"Réunion (NUTS 2010)"
"Y20-64","HU",2001,5.5,"Hungary"
"Y20-64","HU1",2001,4.4,"Közép-Magyarország"
"Y20-64","HU10",2001,4.4,"Közép-Magyarország"
"Y20-64","HU2",2001,4.7,"Dunántúl"
"Y20-64","HU21",2001,3.7,"Közép-Dunántúl"
"Y20-64","HU22",2001,3.6,"Nyugat-Dunántúl"
"Y20-64","HU23",2001,7.2,"Dél-Dunántúl"
"Y20-64","HU3",2001,7,"Alföld és Észak"
"Y20-64","HU31",2001,7.9,"Észak-Magyarország"
"Y20-64","HU32",2001,8.1,"Észak-Alföld"
"Y20-64","HU33",2001,5.3,"Dél-Alföld"
"Y20-64","IE",2001,3.5,"Ireland"
"Y20-64","IE0",2001,3.5,"Éire/Ireland"
"Y20-64","IE01",2001,4.3,"Border, Midland and Western"
"Y20-64","IE02",2001,3.2,"Southern and Eastern"
"Y20-64","IS",2001,1.5,"Iceland"
"Y20-64","IS0",2001,1.5,"Ísland"
"Y20-64","IS00",2001,1.5,"Ísland"
"Y20-64","IT",2001,9.2,"Italy"
"Y20-64","ITC",2001,4.3,"Nord-Ovest"
"Y20-64","ITC1",2001,4.9,"Piemonte"
"Y20-64","ITC2",2001,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2001,5.8,"Liguria"
"Y20-64","ITC4",2001,3.7,"Lombardia"
"Y20-64","ITF",2001,17.4,"Sud"
"Y20-64","ITF1",2001,4.1,"Abruzzo"
"Y20-64","ITF2",2001,12.9,"Molise"
"Y20-64","ITF3",2001,21.5,"Campania"
"Y20-64","ITF4",2001,13.6,"Puglia"
"Y20-64","ITF5",2001,15,"Basilicata"
"Y20-64","ITF6",2001,23.9,"Calabria"
"Y20-64","ITG",2001,19.6,"Isole"
"Y20-64","ITG1",2001,20.1,"Sicilia"
"Y20-64","ITG2",2001,18.4,"Sardegna"
"Y20-64","ITH",2001,3.9,"Nord-Est"
"Y20-64","ITH1",2001,2.2,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2001,3.7,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2001,3.7,"Veneto"
"Y20-64","ITH4",2001,3.7,"Friuli-Venezia Giulia"
"Y20-64","ITI",2001,7.3,"Centro (IT)"
"Y20-64","ITI1",2001,4.8,"Toscana"
"Y20-64","ITI2",2001,4.9,"Umbria"
"Y20-64","ITI4",2001,10.1,"Lazio"
"Y20-64","LT",2001,16.7,"Lithuania"
"Y20-64","LT0",2001,16.7,"Lietuva"
"Y20-64","LT00",2001,16.7,"Lietuva"
"Y20-64","LU",2001,1.7,"Luxembourg"
"Y20-64","LU0",2001,1.7,"Luxembourg"
"Y20-64","LU00",2001,1.7,"Luxembourg"
"Y20-64","LV",2001,13.6,"Latvia"
"Y20-64","LV0",2001,13.6,"Latvija"
"Y20-64","LV00",2001,13.6,"Latvija"
"Y20-64","MT",2001,4.5,"Malta"
"Y20-64","MT0",2001,4.5,"Malta"
"Y20-64","MT00",2001,4.5,"Malta"
"Y20-64","NL",2001,1.8,"Netherlands"
"Y20-64","NL1",2001,2.8,"Noord-Nederland"
"Y20-64","NL11",2001,3.6,"Groningen"
"Y20-64","NL12",2001,2.5,"Friesland (NL)"
"Y20-64","NL13",2001,2.3,"Drenthe"
"Y20-64","NL2",2001,1.9,"Oost-Nederland"
"Y20-64","NL21",2001,2,"Overijssel"
"Y20-64","NL22",2001,1.9,"Gelderland"
"Y20-64","NL23",2001,1.4,"Flevoland"
"Y20-64","NL3",2001,1.6,"West-Nederland"
"Y20-64","NL31",2001,1,"Utrecht"
"Y20-64","NL32",2001,1.7,"Noord-Holland"
"Y20-64","NL33",2001,1.7,"Zuid-Holland"
"Y20-64","NL34",2001,2.6,"Zeeland"
"Y20-64","NL4",2001,1.6,"Zuid-Nederland"
"Y20-64","NL41",2001,1.5,"Noord-Brabant"
"Y20-64","NL42",2001,1.9,"Limburg (NL)"
"Y20-64","NO",2001,2.9,"Norway"
"Y20-64","NO0",2001,2.9,"Norge"
"Y20-64","NO01",2001,2.5,"Oslo og Akershus"
"Y20-64","NO02",2001,2,"Hedmark og Oppland"
"Y20-64","NO03",2001,2.8,"Sør-Østlandet"
"Y20-64","NO04",2001,3.6,"Agder og Rogaland"
"Y20-64","NO05",2001,2.9,"Vestlandet"
"Y20-64","NO06",2001,2.2,"Trøndelag"
"Y20-64","NO07",2001,3.9,"Nord-Norge"
"Y20-64","PL",2001,18.1,"Poland"
"Y20-64","PL1",2001,16.2,"Region Centralny"
"Y20-64","PL11",2001,19.3,"Lódzkie"
"Y20-64","PL12",2001,14.4,"Mazowieckie"
"Y20-64","PL2",2001,16.5,"Region Poludniowy"
"Y20-64","PL21",2001,12.6,"Malopolskie"
"Y20-64","PL22",2001,19.6,"Slaskie"
"Y20-64","PL3",2001,16.5,"Region Wschodni"
"Y20-64","PL31",2001,14.5,"Lubelskie"
"Y20-64","PL32",2001,17.1,"Podkarpackie"
"Y20-64","PL33",2001,19.7,"Swietokrzyskie"
"Y20-64","PL34",2001,16.1,"Podlaskie"
"Y20-64","PL4",2001,19.7,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2001,18.5,"Wielkopolskie"
"Y20-64","PL42",2001,20.5,"Zachodniopomorskie"
"Y20-64","PL43",2001,22.6,"Lubuskie"
"Y20-64","PL5",2001,22.5,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2001,23.9,"Dolnoslaskie"
"Y20-64","PL52",2001,19,"Opolskie"
"Y20-64","PL6",2001,20,"Region Pólnocny"
"Y20-64","PL61",2001,21.5,"Kujawsko-Pomorskie"
"Y20-64","PL62",2001,21.5,"Warminsko-Mazurskie"
"Y20-64","PL63",2001,17.2,"Pomorskie"
"Y20-64","PT",2001,3.8,"Portugal"
"Y20-64","PT1",2001,3.9,"Continente"
"Y20-64","PT11",2001,3.7,"Norte"
"Y20-64","PT15",2001,NA,"Algarve"
"Y20-64","PT16",2001,3,"Centro (PT)"
"Y20-64","PT17",2001,4.7,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2001,5,"Alentejo"
"Y20-64","PT2",2001,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2001,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2001,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2001,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2001,6.9,"Romania"
"Y20-64","RO1",2001,6.6,"Macroregiunea unu"
"Y20-64","RO11",2001,7.2,"Nord-Vest"
"Y20-64","RO12",2001,5.9,"Centru"
"Y20-64","RO2",2001,7.3,"Macroregiunea doi"
"Y20-64","RO21",2001,6.1,"Nord-Est"
"Y20-64","RO22",2001,9,"Sud-Est"
"Y20-64","RO3",2001,7.9,"Macroregiunea trei"
"Y20-64","RO31",2001,7,"Sud - Muntenia"
"Y20-64","RO32",2001,9.3,"Bucuresti - Ilfov"
"Y20-64","RO4",2001,5.3,"Macroregiunea patru"
"Y20-64","RO41",2001,5.5,"Sud-Vest Oltenia"
"Y20-64","RO42",2001,5,"Vest"
"Y20-64","SE",2001,4.2,"Sweden"
"Y20-64","SE1",2001,3.5,"Östra Sverige"
"Y20-64","SE11",2001,2.8,"Stockholm"
"Y20-64","SE12",2001,4.4,"Östra Mellansverige"
"Y20-64","SE2",2001,4.1,"Södra Sverige"
"Y20-64","SE21",2001,3.7,"Småland med öarna"
"Y20-64","SE22",2001,5.3,"Sydsverige"
"Y20-64","SE23",2001,3.6,"Västsverige"
"Y20-64","SE3",2001,6,"Norra Sverige"
"Y20-64","SE31",2001,6,"Norra Mellansverige"
"Y20-64","SE32",2001,6.5,"Mellersta Norrland"
"Y20-64","SE33",2001,5.5,"Övre Norrland"
"Y20-64","SI",2001,5.5,"Slovenia"
"Y20-64","SI0",2001,5.5,"Slovenija"
"Y20-64","SI01",2001,6.4,"Vzhodna Slovenija (NUTS 2010)"
"Y20-64","SI02",2001,4.5,"Zahodna Slovenija (NUTS 2010)"
"Y20-64","SK",2001,18.1,"Slovakia"
"Y20-64","SK0",2001,18.1,"Slovensko"
"Y20-64","SK01",2001,6.8,"Bratislavský kraj"
"Y20-64","SK02",2001,17.2,"Západné Slovensko"
"Y20-64","SK03",2001,20,"Stredné Slovensko"
"Y20-64","SK04",2001,22.7,"Východné Slovensko"
"Y20-64","UK",2001,4.2,"United Kingdom"
"Y20-64","UKC",2001,6.5,"North East (UK)"
"Y20-64","UKC1",2001,6.9,"Tees Valley and Durham"
"Y20-64","UKC2",2001,6.3,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2001,4.2,"North West (UK)"
"Y20-64","UKD1",2001,6,"Cumbria"
"Y20-64","UKD3",2001,3.6,"Greater Manchester"
"Y20-64","UKD4",2001,3.2,"Lancashire"
"Y20-64","UKE",2001,4.2,"Yorkshire and The Humber"
"Y20-64","UKE1",2001,4.7,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2001,NA,"North Yorkshire"
"Y20-64","UKE3",2001,5.3,"South Yorkshire"
"Y20-64","UKE4",2001,4,"West Yorkshire"
"Y20-64","UKF",2001,4.3,"East Midlands (UK)"
"Y20-64","UKF1",2001,4.9,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2001,3.8,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2001,3.9,"Lincolnshire"
"Y20-64","UKG",2001,4.5,"West Midlands (UK)"
"Y20-64","UKG1",2001,2.7,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2001,3.2,"Shropshire and Staffordshire"
"Y20-64","UKG3",2001,6.3,"West Midlands"
"Y20-64","UKH",2001,3,"East of England"
"Y20-64","UKH1",2001,3.3,"East Anglia"
"Y20-64","UKH2",2001,2.6,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2001,3.1,"Essex"
"Y20-64","UKI",2001,5.3,"London"
"Y20-64","UKI1",2001,7.3,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2001,4,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2001,2.6,"South East (UK)"
"Y20-64","UKJ1",2001,2.6,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2001,2.4,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2001,2.1,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2001,3.8,"Kent"
"Y20-64","UKK",2001,3.2,"South West (UK)"
"Y20-64","UKK1",2001,2.7,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2001,2.2,"Dorset and Somerset"
"Y20-64","UKK3",2001,NA,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2001,4.9,"Devon"
"Y20-64","UKL",2001,4.9,"Wales"
"Y20-64","UKL1",2001,5.2,"West Wales and The Valleys"
"Y20-64","UKL2",2001,4.5,"East Wales"
"Y20-64","UKM",2001,4.9,"Scotland"
"Y20-64","UKM2",2001,3.8,"Eastern Scotland"
"Y20-64","UKM3",2001,6.2,"South Western Scotland"
"Y20-64","UKM5",2001,NA,"North Eastern Scotland"
"Y20-64","UKM6",2001,6.5,"Highlands and Islands"
"Y20-64","UKN",2001,5.5,"Northern Ireland (UK)"
"Y20-64","UKN0",2001,5.5,"Northern Ireland (UK)"
"Y_GE15","AT",2001,4,"Austria"
"Y_GE15","AT1",2001,4.7,"Ostösterreich"
"Y_GE15","AT11",2001,5,"Burgenland (AT)"
"Y_GE15","AT12",2001,3.2,"Niederösterreich"
"Y_GE15","AT13",2001,6,"Wien"
"Y_GE15","AT2",2001,4.5,"Südösterreich"
"Y_GE15","AT21",2001,4.6,"Kärnten"
"Y_GE15","AT22",2001,4.5,"Steiermark"
"Y_GE15","AT3",2001,2.9,"Westösterreich"
"Y_GE15","AT31",2001,3.1,"Oberösterreich"
"Y_GE15","AT32",2001,2,"Salzburg"
"Y_GE15","AT33",2001,2.9,"Tirol"
"Y_GE15","AT34",2001,3,"Vorarlberg"
"Y_GE15","BE",2001,6.2,"Belgium"
"Y_GE15","BE1",2001,13,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2001,13,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2001,3.5,"Vlaams Gewest"
"Y_GE15","BE21",2001,4.3,"Prov. Antwerpen"
"Y_GE15","BE22",2001,3.6,"Prov. Limburg (BE)"
"Y_GE15","BE23",2001,3.6,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2001,3.7,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2001,1.9,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2001,9.3,"Région wallonne"
"Y_GE15","BE31",2001,5.9,"Prov. Brabant Wallon"
"Y_GE15","BE32",2001,11.7,"Prov. Hainaut"
"Y_GE15","BE33",2001,9.4,"Prov. Liège"
"Y_GE15","BE34",2001,5.6,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2001,7.8,"Prov. Namur"
"Y_GE15","BG",2001,19.9,"Bulgaria"
"Y_GE15","BG41",2001,15.5,"Yugozapaden"
"Y_GE15","CH",2001,2.5,"Switzerland"
"Y_GE15","CH0",2001,2.5,"Schweiz/Suisse/Svizzera"
"Y_GE15","CH01",2001,4,"Région lémanique"
"Y_GE15","CH02",2001,1.8,"Espace Mittelland"
"Y_GE15","CH03",2001,2.3,"Nordwestschweiz"
"Y_GE15","CH04",2001,2.6,"Zürich"
"Y_GE15","CH05",2001,2,"Ostschweiz"
"Y_GE15","CH06",2001,2.3,"Zentralschweiz"
"Y_GE15","CH07",2001,2.7,"Ticino"
"Y_GE15","CY",2001,4,"Cyprus"
"Y_GE15","CY0",2001,4,"Kypros"
"Y_GE15","CY00",2001,4,"Kypros"
"Y_GE15","CZ",2001,8,"Czech Republic"
"Y_GE15","CZ0",2001,8,"Ceská republika"
"Y_GE15","CZ01",2001,3.8,"Praha"
"Y_GE15","CZ02",2001,6.7,"Strední Cechy"
"Y_GE15","CZ03",2001,5.1,"Jihozápad"
"Y_GE15","CZ04",2001,11.7,"Severozápad"
"Y_GE15","CZ05",2001,5.8,"Severovýchod"
"Y_GE15","CZ06",2001,7.3,"Jihovýchod"
"Y_GE15","CZ07",2001,9.3,"Strední Morava"
"Y_GE15","CZ08",2001,15.2,"Moravskoslezsko"
"Y_GE15","DE",2001,7.8,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2001,3.7,"Baden-Württemberg"
"Y_GE15","DE11",2001,3.6,"Stuttgart"
"Y_GE15","DE12",2001,4.2,"Karlsruhe"
"Y_GE15","DE13",2001,3.7,"Freiburg"
"Y_GE15","DE14",2001,3.4,"Tübingen"
"Y_GE15","DE2",2001,3.8,"Bayern"
"Y_GE15","DE21",2001,2.8,"Oberbayern"
"Y_GE15","DE22",2001,3.8,"Niederbayern"
"Y_GE15","DE23",2001,4.8,"Oberpfalz"
"Y_GE15","DE24",2001,5.4,"Oberfranken"
"Y_GE15","DE25",2001,4.7,"Mittelfranken"
"Y_GE15","DE26",2001,4.3,"Unterfranken"
"Y_GE15","DE27",2001,3.8,"Schwaben"
"Y_GE15","DE3",2001,15.1,"Berlin"
"Y_GE15","DE30",2001,15.1,"Berlin"
"Y_GE15","DE4",2001,16.9,"Brandenburg"
"Y_GE15","DE40",2001,16.9,"Brandenburg"
"Y_GE15","DE5",2001,8.7,"Bremen"
"Y_GE15","DE50",2001,8.7,"Bremen"
"Y_GE15","DE6",2001,7,"Hamburg"
"Y_GE15","DE60",2001,7,"Hamburg"
"Y_GE15","DE7",2001,5.5,"Hessen"
"Y_GE15","DE71",2001,5.1,"Darmstadt"
"Y_GE15","DE72",2001,5.2,"Gießen"
"Y_GE15","DE73",2001,7,"Kassel"
"Y_GE15","DE8",2001,18.5,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2001,18.5,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2001,6.4,"Niedersachsen"
"Y_GE15","DE91",2001,8,"Braunschweig"
"Y_GE15","DE92",2001,6.5,"Hannover"
"Y_GE15","DE93",2001,5.9,"Lüneburg"
"Y_GE15","DE94",2001,5.5,"Weser-Ems"
"Y_GE15","DEA",2001,6,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2001,6,"Düsseldorf"
"Y_GE15","DEA2",2001,5.7,"Köln"
"Y_GE15","DEA3",2001,5.7,"Münster"
"Y_GE15","DEA4",2001,5.7,"Detmold"
"Y_GE15","DEA5",2001,6.9,"Arnsberg"
"Y_GE15","DEB",2001,5,"Rheinland-Pfalz"
"Y_GE15","DEC",2001,5.9,"Saarland"
"Y_GE15","DEC0",2001,5.9,"Saarland"
"Y_GE15","DED",2001,17,"Sachsen"
"Y_GE15","DED2",2001,17.4,"Dresden"
"Y_GE15","DEE",2001,19.9,"Sachsen-Anhalt"
"Y_GE15","DEE0",2001,19.9,"Sachsen-Anhalt"
"Y_GE15","DEF",2001,6.4,"Schleswig-Holstein"
"Y_GE15","DEF0",2001,6.4,"Schleswig-Holstein"
"Y_GE15","DEG",2001,13.9,"Thüringen"
"Y_GE15","DEG0",2001,13.9,"Thüringen"
"Y_GE15","DK",2001,4.2,"Denmark"
"Y_GE15","DK0",2001,4.2,"Danmark"
"Y_GE15","EA17",2001,8.3,"Euro area (17 countries)"
"Y_GE15","EA18",2001,8.3,"Euro area (18 countries)"
"Y_GE15","EA19",2001,8.4,"Euro area (19 countries)"
"Y_GE15","EE",2001,13.1,"Estonia"
"Y_GE15","EE0",2001,13.1,"Eesti"
"Y_GE15","EE00",2001,13.1,"Eesti"
"Y_GE15","EL",2001,10.5,"Greece"
"Y_GE15","EL1",2001,11.3,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2001,9.3,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2001,10.9,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2001,16.2,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2001,12.1,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2001,10.7,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2001,12.6,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2001,7.2,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2001,10.3,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2001,14.1,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2001,8.4,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2001,10.4,"Attiki"
"Y_GE15","EL30",2001,10.4,"Attiki"
"Y_GE15","EL4",2001,7.3,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2001,6.3,"Voreio Aigaio"
"Y_GE15","EL42",2001,9.9,"Notio Aigaio"
"Y_GE15","EL43",2001,6.3,"Kriti"
"Y_GE15","ES",2001,10.3,"Spain"
"Y_GE15","ES1",2001,10.2,"Noroeste (ES)"
"Y_GE15","ES11",2001,11.4,"Galicia"
"Y_GE15","ES12",2001,8.2,"Principado de Asturias"
"Y_GE15","ES13",2001,8,"Cantabria"
"Y_GE15","ES2",2001,7.2,"Noreste (ES)"
"Y_GE15","ES21",2001,9.6,"País Vasco"
"Y_GE15","ES22",2001,4.3,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2001,4.1,"La Rioja"
"Y_GE15","ES24",2001,5,"Aragón"
"Y_GE15","ES3",2001,7.5,"Comunidad de Madrid"
"Y_GE15","ES30",2001,7.5,"Comunidad de Madrid"
"Y_GE15","ES4",2001,10.4,"Centro (ES)"
"Y_GE15","ES41",2001,9.7,"Castilla y León"
"Y_GE15","ES42",2001,9.5,"Castilla-la Mancha"
"Y_GE15","ES43",2001,13.9,"Extremadura"
"Y_GE15","ES5",2001,8.7,"Este (ES)"
"Y_GE15","ES51",2001,8.4,"Cataluña"
"Y_GE15","ES52",2001,9.7,"Comunidad Valenciana"
"Y_GE15","ES53",2001,5.9,"Illes Balears"
"Y_GE15","ES6",2001,16.7,"Sur (ES)"
"Y_GE15","ES61",2001,18.1,"Andalucía"
"Y_GE15","ES62",2001,9.4,"Región de Murcia"
"Y_GE15","ES63",2001,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2001,NA,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2001,10.4,"Canarias (ES)"
"Y_GE15","ES70",2001,10.4,"Canarias (ES)"
"Y_GE15","EU15",2001,7.4,"European Union (15 countries)"
"Y_GE15","EU27",2001,8.6,"European Union (27 countries)"
"Y_GE15","FI",2001,10.3,"Finland"
"Y_GE15","FI1",2001,10.3,"Manner-Suomi"
"Y_GE15","FI19",2001,10.7,"Länsi-Suomi"
"Y_GE15","FI2",2001,NA,"Åland"
"Y_GE15","FI20",2001,NA,"Åland"
"Y_GE15","FR",2001,9.1,"France"
"Y_GE15","FR1",2001,7.4,"Île de France"
"Y_GE15","FR10",2001,7.4,"Île de France"
"Y_GE15","FR2",2001,8.2,"Bassin Parisien"
"Y_GE15","FR21",2001,10,"Champagne-Ardenne"
"Y_GE15","FR22",2001,9.2,"Picardie"
"Y_GE15","FR23",2001,8.9,"Haute-Normandie"
"Y_GE15","FR24",2001,7.3,"Centre (FR)"
"Y_GE15","FR25",2001,7.2,"Basse-Normandie"
"Y_GE15","FR26",2001,6.9,"Bourgogne"
"Y_GE15","FR3",2001,14,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2001,14,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2001,6.6,"Est (FR)"
"Y_GE15","FR41",2001,7.8,"Lorraine"
"Y_GE15","FR42",2001,6.1,"Alsace"
"Y_GE15","FR43",2001,4.9,"Franche-Comté"
"Y_GE15","FR5",2001,7.3,"Ouest (FR)"
"Y_GE15","FR51",2001,7.8,"Pays de la Loire"
"Y_GE15","FR52",2001,6.2,"Bretagne"
"Y_GE15","FR53",2001,8.5,"Poitou-Charentes"
"Y_GE15","FR6",2001,9.4,"Sud-Ouest (FR)"
"Y_GE15","FR61",2001,10.3,"Aquitaine"
"Y_GE15","FR62",2001,8.8,"Midi-Pyrénées"
"Y_GE15","FR63",2001,7.4,"Limousin"
"Y_GE15","FR7",2001,7.2,"Centre-Est (FR)"
"Y_GE15","FR71",2001,7.2,"Rhône-Alpes"
"Y_GE15","FR72",2001,7.5,"Auvergne"
"Y_GE15","FR8",2001,12.8,"Méditerranée"
"Y_GE15","FR81",2001,13.5,"Languedoc-Roussillon"
"Y_GE15","FR82",2001,12.4,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2001,NA,"Corse"
"Y_GE15","FR9",2001,27.8,"Départements d'outre-mer (NUTS 2010)"
"Y_GE15","FR91",2001,25.2,"Guadeloupe (NUTS 2010)"
"Y_GE15","FR92",2001,24,"Martinique (NUTS 2010)"
"Y_GE15","FR93",2001,28.1,"Guyane (NUTS 2010)"
"Y_GE15","FR94",2001,31.5,"Réunion (NUTS 2010)"
"Y_GE15","HU",2001,5.7,"Hungary"
"Y_GE15","HU1",2001,4.5,"Közép-Magyarország"
"Y_GE15","HU10",2001,4.5,"Közép-Magyarország"
"Y_GE15","HU2",2001,4.9,"Dunántúl"
"Y_GE15","HU21",2001,3.9,"Közép-Dunántúl"
"Y_GE15","HU22",2001,3.8,"Nyugat-Dunántúl"
"Y_GE15","HU23",2001,7.5,"Dél-Dunántúl"
"Y_GE15","HU3",2001,7.3,"Alföld és Észak"
"Y_GE15","HU31",2001,8.1,"Észak-Magyarország"
"Y_GE15","HU32",2001,8.3,"Észak-Alföld"
"Y_GE15","HU33",2001,5.5,"Dél-Alföld"
"Y_GE15","IE",2001,3.7,"Ireland"
"Y_GE15","IE0",2001,3.7,"Éire/Ireland"
"Y_GE15","IE01",2001,4.5,"Border, Midland and Western"
"Y_GE15","IE02",2001,3.4,"Southern and Eastern"
"Y_GE15","IS",2001,1.9,"Iceland"
"Y_GE15","IS0",2001,1.9,"Ísland"
"Y_GE15","IS00",2001,1.9,"Ísland"
"Y_GE15","IT",2001,9.6,"Italy"
"Y_GE15","ITC",2001,4.5,"Nord-Ovest"
"Y_GE15","ITC1",2001,5.2,"Piemonte"
"Y_GE15","ITC2",2001,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2001,6.1,"Liguria"
"Y_GE15","ITC4",2001,4,"Lombardia"
"Y_GE15","ITF",2001,18.3,"Sud"
"Y_GE15","ITF1",2001,4.3,"Abruzzo"
"Y_GE15","ITF2",2001,13.2,"Molise"
"Y_GE15","ITF3",2001,22.5,"Campania"
"Y_GE15","ITF4",2001,14.4,"Puglia"
"Y_GE15","ITF5",2001,15.8,"Basilicata"
"Y_GE15","ITF6",2001,25,"Calabria"
"Y_GE15","ITG",2001,20.5,"Isole"
"Y_GE15","ITG1",2001,20.9,"Sicilia"
"Y_GE15","ITG2",2001,19.2,"Sardegna"
"Y_GE15","ITH",2001,4,"Nord-Est"
"Y_GE15","ITH1",2001,2.2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2001,3.9,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2001,3.7,"Veneto"
"Y_GE15","ITH4",2001,3.8,"Friuli-Venezia Giulia"
"Y_GE15","ITI",2001,7.5,"Centro (IT)"
"Y_GE15","ITI1",2001,5,"Toscana"
"Y_GE15","ITI2",2001,4.9,"Umbria"
"Y_GE15","ITI4",2001,10.4,"Lazio"
"Y_GE15","LT",2001,16.8,"Lithuania"
"Y_GE15","LT0",2001,16.8,"Lietuva"
"Y_GE15","LT00",2001,16.8,"Lietuva"
"Y_GE15","LU",2001,1.8,"Luxembourg"
"Y_GE15","LU0",2001,1.8,"Luxembourg"
"Y_GE15","LU00",2001,1.8,"Luxembourg"
"Y_GE15","LV",2001,13.8,"Latvia"
"Y_GE15","LV0",2001,13.8,"Latvija"
"Y_GE15","LV00",2001,13.8,"Latvija"
"Y_GE15","MT",2001,7.1,"Malta"
"Y_GE15","MT0",2001,7.1,"Malta"
"Y_GE15","MT00",2001,7.1,"Malta"
"Y_GE15","NL",2001,2.1,"Netherlands"
"Y_GE15","NL1",2001,3.3,"Noord-Nederland"
"Y_GE15","NL11",2001,3.9,"Groningen"
"Y_GE15","NL12",2001,3.1,"Friesland (NL)"
"Y_GE15","NL13",2001,3,"Drenthe"
"Y_GE15","NL2",2001,2.2,"Oost-Nederland"
"Y_GE15","NL21",2001,2.4,"Overijssel"
"Y_GE15","NL22",2001,2.1,"Gelderland"
"Y_GE15","NL23",2001,1.7,"Flevoland"
"Y_GE15","NL3",2001,1.9,"West-Nederland"
"Y_GE15","NL31",2001,1.2,"Utrecht"
"Y_GE15","NL32",2001,1.9,"Noord-Holland"
"Y_GE15","NL33",2001,2,"Zuid-Holland"
"Y_GE15","NL34",2001,2.5,"Zeeland"
"Y_GE15","NL4",2001,2,"Zuid-Nederland"
"Y_GE15","NL41",2001,1.8,"Noord-Brabant"
"Y_GE15","NL42",2001,2.4,"Limburg (NL)"
"Y_GE15","NO",2001,3.7,"Norway"
"Y_GE15","NO0",2001,3.7,"Norge"
"Y_GE15","NO01",2001,2.9,"Oslo og Akershus"
"Y_GE15","NO02",2001,3,"Hedmark og Oppland"
"Y_GE15","NO03",2001,3.8,"Sør-Østlandet"
"Y_GE15","NO04",2001,4.6,"Agder og Rogaland"
"Y_GE15","NO05",2001,3.6,"Vestlandet"
"Y_GE15","NO06",2001,3.3,"Trøndelag"
"Y_GE15","NO07",2001,5.5,"Nord-Norge"
"Y_GE15","PL",2001,18.4,"Poland"
"Y_GE15","PL1",2001,16.3,"Region Centralny"
"Y_GE15","PL11",2001,19.6,"Lódzkie"
"Y_GE15","PL12",2001,14.3,"Mazowieckie"
"Y_GE15","PL2",2001,17,"Region Poludniowy"
"Y_GE15","PL21",2001,12.9,"Malopolskie"
"Y_GE15","PL22",2001,20.4,"Slaskie"
"Y_GE15","PL3",2001,16.7,"Region Wschodni"
"Y_GE15","PL31",2001,14.7,"Lubelskie"
"Y_GE15","PL32",2001,17.4,"Podkarpackie"
"Y_GE15","PL33",2001,20,"Swietokrzyskie"
"Y_GE15","PL34",2001,15.8,"Podlaskie"
"Y_GE15","PL4",2001,20.4,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2001,18.9,"Wielkopolskie"
"Y_GE15","PL42",2001,21.5,"Zachodniopomorskie"
"Y_GE15","PL43",2001,23.4,"Lubuskie"
"Y_GE15","PL5",2001,22.7,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2001,24.1,"Dolnoslaskie"
"Y_GE15","PL52",2001,19.2,"Opolskie"
"Y_GE15","PL6",2001,20.6,"Region Pólnocny"
"Y_GE15","PL61",2001,21.8,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2001,22.3,"Warminsko-Mazurskie"
"Y_GE15","PL63",2001,17.9,"Pomorskie"
"Y_GE15","PT",2001,3.8,"Portugal"
"Y_GE15","PT1",2001,3.9,"Continente"
"Y_GE15","PT11",2001,3.6,"Norte"
"Y_GE15","PT15",2001,NA,"Algarve"
"Y_GE15","PT16",2001,2.8,"Centro (PT)"
"Y_GE15","PT17",2001,4.9,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2001,5.4,"Alentejo"
"Y_GE15","PT2",2001,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2001,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2001,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2001,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2001,6.6,"Romania"
"Y_GE15","RO1",2001,6.5,"Macroregiunea unu"
"Y_GE15","RO11",2001,6.9,"Nord-Vest"
"Y_GE15","RO12",2001,6,"Centru"
"Y_GE15","RO2",2001,6.8,"Macroregiunea doi"
"Y_GE15","RO21",2001,5.6,"Nord-Est"
"Y_GE15","RO22",2001,8.6,"Sud-Est"
"Y_GE15","RO3",2001,7.6,"Macroregiunea trei"
"Y_GE15","RO31",2001,6.5,"Sud - Muntenia"
"Y_GE15","RO32",2001,9.5,"Bucuresti - Ilfov"
"Y_GE15","RO4",2001,5,"Macroregiunea patru"
"Y_GE15","RO41",2001,5,"Sud-Vest Oltenia"
"Y_GE15","RO42",2001,5,"Vest"
"Y_GE15","SE",2001,4.7,"Sweden"
"Y_GE15","SE1",2001,4,"Östra Sverige"
"Y_GE15","SE11",2001,3.2,"Stockholm"
"Y_GE15","SE12",2001,5.1,"Östra Mellansverige"
"Y_GE15","SE2",2001,4.7,"Södra Sverige"
"Y_GE15","SE21",2001,3.9,"Småland med öarna"
"Y_GE15","SE22",2001,5.9,"Sydsverige"
"Y_GE15","SE23",2001,4.1,"Västsverige"
"Y_GE15","SE3",2001,6.4,"Norra Sverige"
"Y_GE15","SE31",2001,6.6,"Norra Mellansverige"
"Y_GE15","SE32",2001,6.6,"Mellersta Norrland"
"Y_GE15","SE33",2001,6,"Övre Norrland"
"Y_GE15","SI",2001,5.7,"Slovenia"
"Y_GE15","SI0",2001,5.7,"Slovenija"
"Y_GE15","SI01",2001,6.5,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE15","SI02",2001,4.7,"Zahodna Slovenija (NUTS 2010)"
"Y_GE15","SK",2001,19.4,"Slovakia"
"Y_GE15","SK0",2001,19.4,"Slovensko"
"Y_GE15","SK01",2001,7.7,"Bratislavský kraj"
"Y_GE15","SK02",2001,18.6,"Západné Slovensko"
"Y_GE15","SK03",2001,21.1,"Stredné Slovensko"
"Y_GE15","SK04",2001,24.4,"Východné Slovensko"
"Y_GE15","UK",2001,4.7,"United Kingdom"
"Y_GE15","UKC",2001,7.4,"North East (UK)"
"Y_GE15","UKC1",2001,7.4,"Tees Valley and Durham"
"Y_GE15","UKC2",2001,7.4,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2001,5,"North West (UK)"
"Y_GE15","UKD1",2001,6.2,"Cumbria"
"Y_GE15","UKD3",2001,4.1,"Greater Manchester"
"Y_GE15","UKD4",2001,3.7,"Lancashire"
"Y_GE15","UKE",2001,4.7,"Yorkshire and The Humber"
"Y_GE15","UKE1",2001,5.3,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2001,NA,"North Yorkshire"
"Y_GE15","UKE3",2001,5.7,"South Yorkshire"
"Y_GE15","UKE4",2001,4.8,"West Yorkshire"
"Y_GE15","UKF",2001,4.8,"East Midlands (UK)"
"Y_GE15","UKF1",2001,5.5,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2001,4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2001,4.6,"Lincolnshire"
"Y_GE15","UKG",2001,4.9,"West Midlands (UK)"
"Y_GE15","UKG1",2001,2.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2001,3.5,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2001,7,"West Midlands"
"Y_GE15","UKH",2001,3.5,"East of England"
"Y_GE15","UKH1",2001,3.8,"East Anglia"
"Y_GE15","UKH2",2001,3.2,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2001,3.5,"Essex"
"Y_GE15","UKI",2001,5.8,"London"
"Y_GE15","UKI1",2001,7.8,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2001,4.5,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2001,2.9,"South East (UK)"
"Y_GE15","UKJ1",2001,2.9,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2001,2.7,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2001,2.5,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2001,3.9,"Kent"
"Y_GE15","UKK",2001,3.5,"South West (UK)"
"Y_GE15","UKK1",2001,2.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2001,2.6,"Dorset and Somerset"
"Y_GE15","UKK3",2001,4.8,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2001,5,"Devon"
"Y_GE15","UKL",2001,5.5,"Wales"
"Y_GE15","UKL1",2001,5.8,"West Wales and The Valleys"
"Y_GE15","UKL2",2001,5.1,"East Wales"
"Y_GE15","UKM",2001,5.7,"Scotland"
"Y_GE15","UKM2",2001,4.2,"Eastern Scotland"
"Y_GE15","UKM3",2001,7,"South Western Scotland"
"Y_GE15","UKM5",2001,NA,"North Eastern Scotland"
"Y_GE15","UKM6",2001,7.9,"Highlands and Islands"
"Y_GE15","UKN",2001,6.1,"Northern Ireland (UK)"
"Y_GE15","UKN0",2001,6.1,"Northern Ireland (UK)"
"Y_GE25","AT",2001,3.7,"Austria"
"Y_GE25","AT1",2001,4.5,"Ostösterreich"
"Y_GE25","AT11",2001,4.9,"Burgenland (AT)"
"Y_GE25","AT12",2001,2.9,"Niederösterreich"
"Y_GE25","AT13",2001,5.7,"Wien"
"Y_GE25","AT2",2001,3.9,"Südösterreich"
"Y_GE25","AT21",2001,4.1,"Kärnten"
"Y_GE25","AT22",2001,3.8,"Steiermark"
"Y_GE25","AT3",2001,2.7,"Westösterreich"
"Y_GE25","AT31",2001,2.9,"Oberösterreich"
"Y_GE25","AT32",2001,NA,"Salzburg"
"Y_GE25","AT33",2001,2.7,"Tirol"
"Y_GE25","AT34",2001,3.1,"Vorarlberg"
"Y_GE25","BE",2001,5.2,"Belgium"
"Y_GE25","BE1",2001,12.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2001,12.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2001,2.9,"Vlaams Gewest"
"Y_GE25","BE21",2001,3.7,"Prov. Antwerpen"
"Y_GE25","BE22",2001,2.3,"Prov. Limburg (BE)"
"Y_GE25","BE23",2001,3,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2001,3,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2001,2.1,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2001,7.4,"Région wallonne"
"Y_GE25","BE31",2001,4.6,"Prov. Brabant Wallon"
"Y_GE25","BE32",2001,8.8,"Prov. Hainaut"
"Y_GE25","BE33",2001,8,"Prov. Liège"
"Y_GE25","BE34",2001,NA,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2001,6.1,"Prov. Namur"
"Y_GE25","BG",2001,17.6,"Bulgaria"
"Y_GE25","BG41",2001,13.5,"Yugozapaden"
"Y_GE25","CH",2001,2,"Switzerland"
"Y_GE25","CH0",2001,2,"Schweiz/Suisse/Svizzera"
"Y_GE25","CH01",2001,2.8,"Région lémanique"
"Y_GE25","CH02",2001,1.3,"Espace Mittelland"
"Y_GE25","CH03",2001,2.3,"Nordwestschweiz"
"Y_GE25","CH04",2001,2.1,"Zürich"
"Y_GE25","CH05",2001,1.5,"Ostschweiz"
"Y_GE25","CH06",2001,2,"Zentralschweiz"
"Y_GE25","CH07",2001,2.1,"Ticino"
"Y_GE25","CY",2001,3.4,"Cyprus"
"Y_GE25","CY0",2001,3.4,"Kypros"
"Y_GE25","CY00",2001,3.4,"Kypros"
"Y_GE25","CZ",2001,6.9,"Czech Republic"
"Y_GE25","CZ0",2001,6.9,"Ceská republika"
"Y_GE25","CZ01",2001,3.3,"Praha"
"Y_GE25","CZ02",2001,5.8,"Strední Cechy"
"Y_GE25","CZ03",2001,4.8,"Jihozápad"
"Y_GE25","CZ04",2001,10.3,"Severozápad"
"Y_GE25","CZ05",2001,4.7,"Severovýchod"
"Y_GE25","CZ06",2001,6.1,"Jihovýchod"
"Y_GE25","CZ07",2001,8.1,"Strední Morava"
"Y_GE25","CZ08",2001,12.9,"Moravskoslezsko"
"Y_GE25","DE",2001,7.8,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2001,3.7,"Baden-Württemberg"
"Y_GE25","DE11",2001,3.5,"Stuttgart"
"Y_GE25","DE12",2001,4.2,"Karlsruhe"
"Y_GE25","DE13",2001,3.7,"Freiburg"
"Y_GE25","DE14",2001,3.6,"Tübingen"
"Y_GE25","DE2",2001,3.8,"Bayern"
"Y_GE25","DE21",2001,2.7,"Oberbayern"
"Y_GE25","DE22",2001,4,"Niederbayern"
"Y_GE25","DE23",2001,4.9,"Oberpfalz"
"Y_GE25","DE24",2001,5.3,"Oberfranken"
"Y_GE25","DE25",2001,4.7,"Mittelfranken"
"Y_GE25","DE26",2001,4.4,"Unterfranken"
"Y_GE25","DE27",2001,3.7,"Schwaben"
"Y_GE25","DE3",2001,14.8,"Berlin"
"Y_GE25","DE30",2001,14.8,"Berlin"
"Y_GE25","DE4",2001,17.3,"Brandenburg"
"Y_GE25","DE40",2001,17.3,"Brandenburg"
"Y_GE25","DE5",2001,8.5,"Bremen"
"Y_GE25","DE50",2001,8.5,"Bremen"
"Y_GE25","DE6",2001,6.8,"Hamburg"
"Y_GE25","DE60",2001,6.8,"Hamburg"
"Y_GE25","DE7",2001,5.5,"Hessen"
"Y_GE25","DE71",2001,5.1,"Darmstadt"
"Y_GE25","DE72",2001,5.2,"Gießen"
"Y_GE25","DE73",2001,6.8,"Kassel"
"Y_GE25","DE8",2001,19.5,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2001,19.5,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2001,6.2,"Niedersachsen"
"Y_GE25","DE91",2001,7.7,"Braunschweig"
"Y_GE25","DE92",2001,6.7,"Hannover"
"Y_GE25","DE93",2001,5.4,"Lüneburg"
"Y_GE25","DE94",2001,5.2,"Weser-Ems"
"Y_GE25","DEA",2001,6,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2001,5.9,"Düsseldorf"
"Y_GE25","DEA2",2001,5.5,"Köln"
"Y_GE25","DEA3",2001,5.7,"Münster"
"Y_GE25","DEA4",2001,5.8,"Detmold"
"Y_GE25","DEA5",2001,6.7,"Arnsberg"
"Y_GE25","DEB",2001,4.8,"Rheinland-Pfalz"
"Y_GE25","DEC",2001,6,"Saarland"
"Y_GE25","DEC0",2001,6,"Saarland"
"Y_GE25","DED",2001,17.5,"Sachsen"
"Y_GE25","DED2",2001,17.5,"Dresden"
"Y_GE25","DEE",2001,20.8,"Sachsen-Anhalt"
"Y_GE25","DEE0",2001,20.8,"Sachsen-Anhalt"
"Y_GE25","DEF",2001,6.1,"Schleswig-Holstein"
"Y_GE25","DEF0",2001,6.1,"Schleswig-Holstein"
"Y_GE25","DEG",2001,14.2,"Thüringen"
"Y_GE25","DEG0",2001,14.2,"Thüringen"
"Y_GE25","DK",2001,3.5,"Denmark"
"Y_GE25","DK0",2001,3.5,"Danmark"
"Y_GE25","EA17",2001,7.3,"Euro area (17 countries)"
"Y_GE25","EA18",2001,7.3,"Euro area (18 countries)"
"Y_GE25","EA19",2001,7.4,"Euro area (19 countries)"
"Y_GE25","EE",2001,11.9,"Estonia"
"Y_GE25","EE0",2001,11.9,"Eesti"
"Y_GE25","EE00",2001,11.9,"Eesti"
"Y_GE25","EL",2001,8.2,"Greece"
"Y_GE25","EL1",2001,9.2,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2001,7.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2001,8.6,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2001,13.5,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2001,10,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2001,8,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2001,10.1,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2001,6.2,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2001,7,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2001,10.1,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2001,6.6,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2001,8.3,"Attiki"
"Y_GE25","EL30",2001,8.3,"Attiki"
"Y_GE25","EL4",2001,5.4,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2001,4.4,"Voreio Aigaio"
"Y_GE25","EL42",2001,8.2,"Notio Aigaio"
"Y_GE25","EL43",2001,4.4,"Kriti"
"Y_GE25","ES",2001,8.7,"Spain"
"Y_GE25","ES1",2001,8.7,"Noroeste (ES)"
"Y_GE25","ES11",2001,9.5,"Galicia"
"Y_GE25","ES12",2001,7.3,"Principado de Asturias"
"Y_GE25","ES13",2001,7.5,"Cantabria"
"Y_GE25","ES2",2001,6.2,"Noreste (ES)"
"Y_GE25","ES21",2001,8.1,"País Vasco"
"Y_GE25","ES22",2001,3.5,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2001,3.4,"La Rioja"
"Y_GE25","ES24",2001,4.4,"Aragón"
"Y_GE25","ES3",2001,6.1,"Comunidad de Madrid"
"Y_GE25","ES30",2001,6.1,"Comunidad de Madrid"
"Y_GE25","ES4",2001,8.8,"Centro (ES)"
"Y_GE25","ES41",2001,8,"Castilla y León"
"Y_GE25","ES42",2001,7.8,"Castilla-la Mancha"
"Y_GE25","ES43",2001,12.6,"Extremadura"
"Y_GE25","ES5",2001,7.3,"Este (ES)"
"Y_GE25","ES51",2001,7.2,"Cataluña"
"Y_GE25","ES52",2001,8.2,"Comunidad Valenciana"
"Y_GE25","ES53",2001,4.5,"Illes Balears"
"Y_GE25","ES6",2001,14.4,"Sur (ES)"
"Y_GE25","ES61",2001,15.7,"Andalucía"
"Y_GE25","ES62",2001,7.5,"Región de Murcia"
"Y_GE25","ES63",2001,NA,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2001,NA,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2001,8.7,"Canarias (ES)"
"Y_GE25","ES70",2001,8.7,"Canarias (ES)"
"Y_GE25","EU15",2001,6.4,"European Union (15 countries)"
"Y_GE25","EU27",2001,7.4,"European Union (27 countries)"
"Y_GE25","FI",2001,7.4,"Finland"
"Y_GE25","FI1",2001,7.5,"Manner-Suomi"
"Y_GE25","FI19",2001,7.4,"Länsi-Suomi"
"Y_GE25","FI2",2001,NA,"Åland"
"Y_GE25","FI20",2001,NA,"Åland"
"Y_GE25","FR",2001,8,"France"
"Y_GE25","FR1",2001,6.7,"Île de France"
"Y_GE25","FR10",2001,6.7,"Île de France"
"Y_GE25","FR2",2001,7.1,"Bassin Parisien"
"Y_GE25","FR21",2001,8.6,"Champagne-Ardenne"
"Y_GE25","FR22",2001,7.7,"Picardie"
"Y_GE25","FR23",2001,7.7,"Haute-Normandie"
"Y_GE25","FR24",2001,6.3,"Centre (FR)"
"Y_GE25","FR25",2001,6.2,"Basse-Normandie"
"Y_GE25","FR26",2001,6.5,"Bourgogne"
"Y_GE25","FR3",2001,12.1,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2001,12.1,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2001,5.7,"Est (FR)"
"Y_GE25","FR41",2001,6.8,"Lorraine"
"Y_GE25","FR42",2001,5,"Alsace"
"Y_GE25","FR43",2001,4.3,"Franche-Comté"
"Y_GE25","FR5",2001,6.5,"Ouest (FR)"
"Y_GE25","FR51",2001,6.9,"Pays de la Loire"
"Y_GE25","FR52",2001,5.5,"Bretagne"
"Y_GE25","FR53",2001,8,"Poitou-Charentes"
"Y_GE25","FR6",2001,8.1,"Sud-Ouest (FR)"
"Y_GE25","FR61",2001,8.9,"Aquitaine"
"Y_GE25","FR62",2001,7.5,"Midi-Pyrénées"
"Y_GE25","FR63",2001,6.2,"Limousin"
"Y_GE25","FR7",2001,6.3,"Centre-Est (FR)"
"Y_GE25","FR71",2001,6.3,"Rhône-Alpes"
"Y_GE25","FR72",2001,6.3,"Auvergne"
"Y_GE25","FR8",2001,11.3,"Méditerranée"
"Y_GE25","FR81",2001,11.5,"Languedoc-Roussillon"
"Y_GE25","FR82",2001,11.2,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2001,NA,"Corse"
"Y_GE25","FR9",2001,24.6,"Départements d'outre-mer (NUTS 2010)"
"Y_GE25","FR91",2001,22.6,"Guadeloupe (NUTS 2010)"
"Y_GE25","FR92",2001,21.6,"Martinique (NUTS 2010)"
"Y_GE25","FR93",2001,25.4,"Guyane (NUTS 2010)"
"Y_GE25","FR94",2001,27.6,"Réunion (NUTS 2010)"
"Y_GE25","HU",2001,5,"Hungary"
"Y_GE25","HU1",2001,3.9,"Közép-Magyarország"
"Y_GE25","HU10",2001,3.9,"Közép-Magyarország"
"Y_GE25","HU2",2001,4.3,"Dunántúl"
"Y_GE25","HU21",2001,3.7,"Közép-Dunántúl"
"Y_GE25","HU22",2001,3.1,"Nyugat-Dunántúl"
"Y_GE25","HU23",2001,6.5,"Dél-Dunántúl"
"Y_GE25","HU3",2001,6.5,"Alföld és Észak"
"Y_GE25","HU31",2001,7.3,"Észak-Magyarország"
"Y_GE25","HU32",2001,7.5,"Észak-Alföld"
"Y_GE25","HU33",2001,4.7,"Dél-Alföld"
"Y_GE25","IE",2001,3.1,"Ireland"
"Y_GE25","IE0",2001,3.1,"Éire/Ireland"
"Y_GE25","IE01",2001,3.9,"Border, Midland and Western"
"Y_GE25","IE02",2001,2.9,"Southern and Eastern"
"Y_GE25","IS",2001,1.2,"Iceland"
"Y_GE25","IS0",2001,1.2,"Ísland"
"Y_GE25","IS00",2001,1.2,"Ísland"
"Y_GE25","IT",2001,7.6,"Italy"
"Y_GE25","ITC",2001,3.6,"Nord-Ovest"
"Y_GE25","ITC1",2001,4.3,"Piemonte"
"Y_GE25","ITC2",2001,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2001,4.6,"Liguria"
"Y_GE25","ITC4",2001,3.2,"Lombardia"
"Y_GE25","ITF",2001,14.1,"Sud"
"Y_GE25","ITF1",2001,3.1,"Abruzzo"
"Y_GE25","ITF2",2001,10.5,"Molise"
"Y_GE25","ITF3",2001,17.2,"Campania"
"Y_GE25","ITF4",2001,10.9,"Puglia"
"Y_GE25","ITF5",2001,12.6,"Basilicata"
"Y_GE25","ITF6",2001,20.4,"Calabria"
"Y_GE25","ITG",2001,16.3,"Isole"
"Y_GE25","ITG1",2001,16.8,"Sicilia"
"Y_GE25","ITG2",2001,14.8,"Sardegna"
"Y_GE25","ITH",2001,3.5,"Nord-Est"
"Y_GE25","ITH1",2001,1.9,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2001,3.5,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2001,3.3,"Veneto"
"Y_GE25","ITH4",2001,3.5,"Friuli-Venezia Giulia"
"Y_GE25","ITI",2001,6,"Centro (IT)"
"Y_GE25","ITI1",2001,3.9,"Toscana"
"Y_GE25","ITI2",2001,4.2,"Umbria"
"Y_GE25","ITI4",2001,8.4,"Lazio"
"Y_GE25","LT",2001,15.2,"Lithuania"
"Y_GE25","LT0",2001,15.2,"Lietuva"
"Y_GE25","LT00",2001,15.2,"Lietuva"
"Y_GE25","LU",2001,1.3,"Luxembourg"
"Y_GE25","LU0",2001,1.3,"Luxembourg"
"Y_GE25","LU00",2001,1.3,"Luxembourg"
"Y_GE25","LV",2001,12.5,"Latvia"
"Y_GE25","LV0",2001,12.5,"Latvija"
"Y_GE25","LV00",2001,12.5,"Latvija"
"Y_GE25","MT",2001,3.8,"Malta"
"Y_GE25","MT0",2001,3.8,"Malta"
"Y_GE25","MT00",2001,3.8,"Malta"
"Y_GE25","NL",2001,1.7,"Netherlands"
"Y_GE25","NL1",2001,2.6,"Noord-Nederland"
"Y_GE25","NL11",2001,3.1,"Groningen"
"Y_GE25","NL12",2001,2.2,"Friesland (NL)"
"Y_GE25","NL13",2001,2.3,"Drenthe"
"Y_GE25","NL2",2001,1.8,"Oost-Nederland"
"Y_GE25","NL21",2001,1.7,"Overijssel"
"Y_GE25","NL22",2001,1.8,"Gelderland"
"Y_GE25","NL23",2001,1.4,"Flevoland"
"Y_GE25","NL3",2001,1.5,"West-Nederland"
"Y_GE25","NL31",2001,1,"Utrecht"
"Y_GE25","NL32",2001,1.4,"Noord-Holland"
"Y_GE25","NL33",2001,1.6,"Zuid-Holland"
"Y_GE25","NL34",2001,2.6,"Zeeland"
"Y_GE25","NL4",2001,1.5,"Zuid-Nederland"
"Y_GE25","NL41",2001,1.4,"Noord-Brabant"
"Y_GE25","NL42",2001,1.8,"Limburg (NL)"
"Y_GE25","NO",2001,2.3,"Norway"
"Y_GE25","NO0",2001,2.3,"Norge"
"Y_GE25","NO01",2001,2.3,"Oslo og Akershus"
"Y_GE25","NO02",2001,1.4,"Hedmark og Oppland"
"Y_GE25","NO03",2001,2.5,"Sør-Østlandet"
"Y_GE25","NO04",2001,2.9,"Agder og Rogaland"
"Y_GE25","NO05",2001,2.2,"Vestlandet"
"Y_GE25","NO06",2001,1.9,"Trøndelag"
"Y_GE25","NO07",2001,2.8,"Nord-Norge"
"Y_GE25","PL",2001,15.1,"Poland"
"Y_GE25","PL1",2001,13.6,"Region Centralny"
"Y_GE25","PL11",2001,16.4,"Lódzkie"
"Y_GE25","PL12",2001,11.9,"Mazowieckie"
"Y_GE25","PL2",2001,13.6,"Region Poludniowy"
"Y_GE25","PL21",2001,9.4,"Malopolskie"
"Y_GE25","PL22",2001,17,"Slaskie"
"Y_GE25","PL3",2001,13,"Region Wschodni"
"Y_GE25","PL31",2001,11.3,"Lubelskie"
"Y_GE25","PL32",2001,13.2,"Podkarpackie"
"Y_GE25","PL33",2001,15.6,"Swietokrzyskie"
"Y_GE25","PL34",2001,13,"Podlaskie"
"Y_GE25","PL4",2001,16.8,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2001,15.3,"Wielkopolskie"
"Y_GE25","PL42",2001,18,"Zachodniopomorskie"
"Y_GE25","PL43",2001,19.8,"Lubuskie"
"Y_GE25","PL5",2001,19.3,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2001,21,"Dolnoslaskie"
"Y_GE25","PL52",2001,15.4,"Opolskie"
"Y_GE25","PL6",2001,17.5,"Region Pólnocny"
"Y_GE25","PL61",2001,18.9,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2001,18.3,"Warminsko-Mazurskie"
"Y_GE25","PL63",2001,15.1,"Pomorskie"
"Y_GE25","PT",2001,3.1,"Portugal"
"Y_GE25","PT1",2001,3.1,"Continente"
"Y_GE25","PT11",2001,3.2,"Norte"
"Y_GE25","PT15",2001,NA,"Algarve"
"Y_GE25","PT16",2001,2,"Centro (PT)"
"Y_GE25","PT17",2001,3.9,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2001,4.1,"Alentejo"
"Y_GE25","PT2",2001,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2001,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2001,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2001,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2001,5,"Romania"
"Y_GE25","RO1",2001,5.2,"Macroregiunea unu"
"Y_GE25","RO11",2001,6,"Nord-Vest"
"Y_GE25","RO12",2001,4.4,"Centru"
"Y_GE25","RO2",2001,5.1,"Macroregiunea doi"
"Y_GE25","RO21",2001,4.1,"Nord-Est"
"Y_GE25","RO22",2001,6.6,"Sud-Est"
"Y_GE25","RO3",2001,5.7,"Macroregiunea trei"
"Y_GE25","RO31",2001,4.4,"Sud - Muntenia"
"Y_GE25","RO32",2001,8.1,"Bucuresti - Ilfov"
"Y_GE25","RO4",2001,3.9,"Macroregiunea patru"
"Y_GE25","RO41",2001,3.6,"Sud-Vest Oltenia"
"Y_GE25","RO42",2001,4.3,"Vest"
"Y_GE25","SE",2001,3.8,"Sweden"
"Y_GE25","SE1",2001,3.1,"Östra Sverige"
"Y_GE25","SE11",2001,2.4,"Stockholm"
"Y_GE25","SE12",2001,3.9,"Östra Mellansverige"
"Y_GE25","SE2",2001,3.7,"Södra Sverige"
"Y_GE25","SE21",2001,3.3,"Småland med öarna"
"Y_GE25","SE22",2001,4.8,"Sydsverige"
"Y_GE25","SE23",2001,3.2,"Västsverige"
"Y_GE25","SE3",2001,5.5,"Norra Sverige"
"Y_GE25","SE31",2001,5.5,"Norra Mellansverige"
"Y_GE25","SE32",2001,6.1,"Mellersta Norrland"
"Y_GE25","SE33",2001,5.2,"Övre Norrland"
"Y_GE25","SI",2001,4.5,"Slovenia"
"Y_GE25","SI0",2001,4.5,"Slovenija"
"Y_GE25","SI01",2001,5.2,"Vzhodna Slovenija (NUTS 2010)"
"Y_GE25","SI02",2001,3.7,"Zahodna Slovenija (NUTS 2010)"
"Y_GE25","SK",2001,15.8,"Slovakia"
"Y_GE25","SK0",2001,15.8,"Slovensko"
"Y_GE25","SK01",2001,5.7,"Bratislavský kraj"
"Y_GE25","SK02",2001,15.4,"Západné Slovensko"
"Y_GE25","SK03",2001,17.5,"Stredné Slovensko"
"Y_GE25","SK04",2001,19.7,"Východné Slovensko"
"Y_GE25","UK",2001,3.7,"United Kingdom"
"Y_GE25","UKC",2001,6.1,"North East (UK)"
"Y_GE25","UKC1",2001,6.5,"Tees Valley and Durham"
"Y_GE25","UKC2",2001,5.8,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2001,3.6,"North West (UK)"
"Y_GE25","UKD1",2001,NA,"Cumbria"
"Y_GE25","UKD3",2001,2.8,"Greater Manchester"
"Y_GE25","UKD4",2001,2.9,"Lancashire"
"Y_GE25","UKE",2001,3.8,"Yorkshire and The Humber"
"Y_GE25","UKE1",2001,4.3,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2001,NA,"North Yorkshire"
"Y_GE25","UKE3",2001,4.8,"South Yorkshire"
"Y_GE25","UKE4",2001,3.6,"West Yorkshire"
"Y_GE25","UKF",2001,3.8,"East Midlands (UK)"
"Y_GE25","UKF1",2001,4.2,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2001,3.3,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2001,3.8,"Lincolnshire"
"Y_GE25","UKG",2001,4.1,"West Midlands (UK)"
"Y_GE25","UKG1",2001,2.4,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2001,3,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2001,5.8,"West Midlands"
"Y_GE25","UKH",2001,2.7,"East of England"
"Y_GE25","UKH1",2001,2.7,"East Anglia"
"Y_GE25","UKH2",2001,2.5,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2001,3,"Essex"
"Y_GE25","UKI",2001,4.8,"London"
"Y_GE25","UKI1",2001,6.5,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2001,3.6,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2001,2.3,"South East (UK)"
"Y_GE25","UKJ1",2001,2.3,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2001,2.1,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2001,2,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2001,3.1,"Kent"
"Y_GE25","UKK",2001,2.9,"South West (UK)"
"Y_GE25","UKK1",2001,2.6,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2001,NA,"Dorset and Somerset"
"Y_GE25","UKK3",2001,NA,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2001,4.2,"Devon"
"Y_GE25","UKL",2001,4,"Wales"
"Y_GE25","UKL1",2001,4,"West Wales and The Valleys"
"Y_GE25","UKL2",2001,4.1,"East Wales"
"Y_GE25","UKM",2001,4.3,"Scotland"
"Y_GE25","UKM2",2001,2.9,"Eastern Scotland"
"Y_GE25","UKM3",2001,5.7,"South Western Scotland"
"Y_GE25","UKM5",2001,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2001,6.3,"Highlands and Islands"
"Y_GE25","UKN",2001,5.4,"Northern Ireland (UK)"
"Y_GE25","UKN0",2001,5.4,"Northern Ireland (UK)"
"Y15-24","AT",2000,6.3,"Austria"
"Y15-24","AT1",2000,6.6,"Ostösterreich"
"Y15-24","AT11",2000,NA,"Burgenland (AT)"
"Y15-24","AT12",2000,4.4,"Niederösterreich"
"Y15-24","AT13",2000,9.5,"Wien"
"Y15-24","AT2",2000,8,"Südösterreich"
"Y15-24","AT21",2000,NA,"Kärnten"
"Y15-24","AT22",2000,8.4,"Steiermark"
"Y15-24","AT3",2000,5.2,"Westösterreich"
"Y15-24","AT31",2000,6,"Oberösterreich"
"Y15-24","AT32",2000,NA,"Salzburg"
"Y15-24","AT33",2000,NA,"Tirol"
"Y15-24","AT34",2000,NA,"Vorarlberg"
"Y15-24","BE",2000,15.2,"Belgium"
"Y15-24","BE1",2000,34.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",2000,34.4,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",2000,9,"Vlaams Gewest"
"Y15-24","BE21",2000,10.7,"Prov. Antwerpen"
"Y15-24","BE22",2000,NA,"Prov. Limburg (BE)"
"Y15-24","BE23",2000,NA,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",2000,NA,"Prov. Vlaams-Brabant"
"Y15-24","BE25",2000,NA,"Prov. West-Vlaanderen"
"Y15-24","BE3",2000,22.8,"Région wallonne"
"Y15-24","BE31",2000,NA,"Prov. Brabant Wallon"
"Y15-24","BE32",2000,29.6,"Prov. Hainaut"
"Y15-24","BE33",2000,14,"Prov. Liège"
"Y15-24","BE34",2000,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",2000,27,"Prov. Namur"
"Y15-24","BG",2000,33.3,"Bulgaria"
"Y15-24","BG41",2000,23.3,"Yugozapaden"
"Y15-24","CH",2000,5,"Switzerland"
"Y15-24","CH0",2000,5,"Schweiz/Suisse/Svizzera"
"Y15-24","CY",2000,10.2,"Cyprus"
"Y15-24","CY0",2000,10.2,"Kypros"
"Y15-24","CY00",2000,10.2,"Kypros"
"Y15-24","CZ",2000,17,"Czech Republic"
"Y15-24","CZ0",2000,17,"Ceská republika"
"Y15-24","CZ01",2000,11.3,"Praha"
"Y15-24","CZ02",2000,11.6,"Strední Cechy"
"Y15-24","CZ03",2000,10.8,"Jihozápad"
"Y15-24","CZ04",2000,25.6,"Severozápad"
"Y15-24","CZ05",2000,14.3,"Severovýchod"
"Y15-24","CZ06",2000,12.7,"Jihovýchod"
"Y15-24","CZ07",2000,20,"Strední Morava"
"Y15-24","CZ08",2000,30.5,"Moravskoslezsko"
"Y15-24","DE",2000,8.5,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",2000,5.7,"Baden-Württemberg"
"Y15-24","DE11",2000,4.9,"Stuttgart"
"Y15-24","DE12",2000,7.1,"Karlsruhe"
"Y15-24","DE13",2000,7.1,"Freiburg"
"Y15-24","DE14",2000,NA,"Tübingen"
"Y15-24","DE2",2000,4.6,"Bayern"
"Y15-24","DE21",2000,4,"Oberbayern"
"Y15-24","DE22",2000,NA,"Niederbayern"
"Y15-24","DE23",2000,NA,"Oberpfalz"
"Y15-24","DE24",2000,7.2,"Oberfranken"
"Y15-24","DE25",2000,5.3,"Mittelfranken"
"Y15-24","DE26",2000,6.3,"Unterfranken"
"Y15-24","DE27",2000,NA,"Schwaben"
"Y15-24","DE3",2000,15.5,"Berlin"
"Y15-24","DE30",2000,15.5,"Berlin"
"Y15-24","DE4",2000,18.5,"Brandenburg"
"Y15-24","DE40",2000,18.5,"Brandenburg"
"Y15-24","DE5",2000,NA,"Bremen"
"Y15-24","DE50",2000,NA,"Bremen"
"Y15-24","DE6",2000,8.7,"Hamburg"
"Y15-24","DE60",2000,8.7,"Hamburg"
"Y15-24","DE7",2000,6.8,"Hessen"
"Y15-24","DE71",2000,6.1,"Darmstadt"
"Y15-24","DE72",2000,9.3,"Gießen"
"Y15-24","DE73",2000,NA,"Kassel"
"Y15-24","DE8",2000,12,"Mecklenburg-Vorpommern"
"Y15-24","DE80",2000,12,"Mecklenburg-Vorpommern"
"Y15-24","DE9",2000,9.4,"Niedersachsen"
"Y15-24","DE91",2000,11.5,"Braunschweig"
"Y15-24","DE92",2000,9.5,"Hannover"
"Y15-24","DE93",2000,9.1,"Lüneburg"
"Y15-24","DE94",2000,8.2,"Weser-Ems"
"Y15-24","DEA",2000,8,"Nordrhein-Westfalen"
"Y15-24","DEA1",2000,9.5,"Düsseldorf"
"Y15-24","DEA2",2000,7.4,"Köln"
"Y15-24","DEA3",2000,5.5,"Münster"
"Y15-24","DEA4",2000,6.8,"Detmold"
"Y15-24","DEA5",2000,9.5,"Arnsberg"
"Y15-24","DEB",2000,8,"Rheinland-Pfalz"
"Y15-24","DEC",2000,10.6,"Saarland"
"Y15-24","DEC0",2000,10.6,"Saarland"
"Y15-24","DED",2000,12.7,"Sachsen"
"Y15-24","DED2",2000,11.7,"Dresden"
"Y15-24","DEE",2000,12.7,"Sachsen-Anhalt"
"Y15-24","DEE0",2000,12.7,"Sachsen-Anhalt"
"Y15-24","DEF",2000,7.1,"Schleswig-Holstein"
"Y15-24","DEF0",2000,7.1,"Schleswig-Holstein"
"Y15-24","DEG",2000,10.2,"Thüringen"
"Y15-24","DEG0",2000,10.2,"Thüringen"
"Y15-24","DK",2000,6.7,"Denmark"
"Y15-24","DK0",2000,6.7,"Danmark"
"Y15-24","EA17",2000,18,"Euro area (17 countries)"
"Y15-24","EA18",2000,18,"Euro area (18 countries)"
"Y15-24","EA19",2000,18.1,"Euro area (19 countries)"
"Y15-24","EE",2000,21.1,"Estonia"
"Y15-24","EE0",2000,21.1,"Eesti"
"Y15-24","EE00",2000,21.1,"Eesti"
"Y15-24","EL",2000,29.2,"Greece"
"Y15-24","EL1",2000,28.6,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",2000,19.3,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",2000,28.7,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",2000,45.2,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",2000,31.6,"Thessalia (NUTS 2010)"
"Y15-24","EL2",2000,32.7,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",2000,29.9,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",2000,NA,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",2000,34.1,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",2000,41.2,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",2000,29.6,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",2000,30.4,"Attiki"
"Y15-24","EL30",2000,30.4,"Attiki"
"Y15-24","EL4",2000,21,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",2000,NA,"Voreio Aigaio"
"Y15-24","EL42",2000,21.4,"Notio Aigaio"
"Y15-24","EL43",2000,21.6,"Kriti"
"Y15-24","ES",2000,25.3,"Spain"
"Y15-24","ES1",2000,29.8,"Noroeste (ES)"
"Y15-24","ES11",2000,28.1,"Galicia"
"Y15-24","ES12",2000,34.4,"Principado de Asturias"
"Y15-24","ES13",2000,30.8,"Cantabria"
"Y15-24","ES2",2000,20.1,"Noreste (ES)"
"Y15-24","ES21",2000,24.5,"País Vasco"
"Y15-24","ES22",2000,13.2,"Comunidad Foral de Navarra"
"Y15-24","ES23",2000,19.1,"La Rioja"
"Y15-24","ES24",2000,16.6,"Aragón"
"Y15-24","ES3",2000,23.1,"Comunidad de Madrid"
"Y15-24","ES30",2000,23.1,"Comunidad de Madrid"
"Y15-24","ES4",2000,26.9,"Centro (ES)"
"Y15-24","ES41",2000,29.7,"Castilla y León"
"Y15-24","ES42",2000,19.6,"Castilla-la Mancha"
"Y15-24","ES43",2000,33.8,"Extremadura"
"Y15-24","ES5",2000,18.7,"Este (ES)"
"Y15-24","ES51",2000,18.7,"Cataluña"
"Y15-24","ES52",2000,20.6,"Comunidad Valenciana"
"Y15-24","ES53",2000,10,"Illes Balears"
"Y15-24","ES6",2000,34.3,"Sur (ES)"
"Y15-24","ES61",2000,36.4,"Andalucía"
"Y15-24","ES62",2000,22.2,"Región de Murcia"
"Y15-24","ES63",2000,46.5,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",2000,NA,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",2000,24.3,"Canarias (ES)"
"Y15-24","ES70",2000,24.3,"Canarias (ES)"
"Y15-24","EU15",2000,16.1,"European Union (15 countries)"
"Y15-24","EU27",2000,18.3,"European Union (27 countries)"
"Y15-24","FI",2000,28.4,"Finland"
"Y15-24","FI1",2000,28.4,"Manner-Suomi"
"Y15-24","FI19",2000,29.1,"Länsi-Suomi"
"Y15-24","FI2",2000,NA,"Åland"
"Y15-24","FI20",2000,NA,"Åland"
"Y15-24","FR",2000,20.6,"France"
"Y15-24","FR1",2000,16,"Île de France"
"Y15-24","FR10",2000,16,"Île de France"
"Y15-24","FR2",2000,19.9,"Bassin Parisien"
"Y15-24","FR21",2000,24.9,"Champagne-Ardenne"
"Y15-24","FR22",2000,25.6,"Picardie"
"Y15-24","FR23",2000,19.8,"Haute-Normandie"
"Y15-24","FR24",2000,16.7,"Centre (FR)"
"Y15-24","FR25",2000,NA,"Basse-Normandie"
"Y15-24","FR26",2000,16.4,"Bourgogne"
"Y15-24","FR3",2000,37.9,"Nord - Pas-de-Calais"
"Y15-24","FR30",2000,37.9,"Nord - Pas-de-Calais"
"Y15-24","FR4",2000,16.2,"Est (FR)"
"Y15-24","FR41",2000,19.1,"Lorraine"
"Y15-24","FR42",2000,12.2,"Alsace"
"Y15-24","FR43",2000,NA,"Franche-Comté"
"Y15-24","FR5",2000,17.1,"Ouest (FR)"
"Y15-24","FR51",2000,16.2,"Pays de la Loire"
"Y15-24","FR52",2000,18.2,"Bretagne"
"Y15-24","FR53",2000,17.7,"Poitou-Charentes"
"Y15-24","FR6",2000,22.4,"Sud-Ouest (FR)"
"Y15-24","FR61",2000,25.2,"Aquitaine"
"Y15-24","FR62",2000,20.8,"Midi-Pyrénées"
"Y15-24","FR63",2000,NA,"Limousin"
"Y15-24","FR7",2000,17.8,"Centre-Est (FR)"
"Y15-24","FR71",2000,16.6,"Rhône-Alpes"
"Y15-24","FR72",2000,23.6,"Auvergne"
"Y15-24","FR8",2000,26.3,"Méditerranée"
"Y15-24","FR81",2000,34.2,"Languedoc-Roussillon"
"Y15-24","FR82",2000,20.5,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",2000,NA,"Corse"
"Y15-24","HU",2000,12.3,"Hungary"
"Y15-24","HU1",2000,11.6,"Közép-Magyarország"
"Y15-24","HU10",2000,11.6,"Közép-Magyarország"
"Y15-24","HU2",2000,9.4,"Dunántúl"
"Y15-24","HU21",2000,8,"Közép-Dunántúl"
"Y15-24","HU22",2000,8.4,"Nyugat-Dunántúl"
"Y15-24","HU23",2000,12.4,"Dél-Dunántúl"
"Y15-24","HU3",2000,15.1,"Alföld és Észak"
"Y15-24","HU31",2000,20.2,"Észak-Magyarország"
"Y15-24","HU32",2000,16.7,"Észak-Alföld"
"Y15-24","HU33",2000,8,"Dél-Alföld"
"Y15-24","IE",2000,6.5,"Ireland"
"Y15-24","IE0",2000,6.5,"Éire/Ireland"
"Y15-24","IE01",2000,9.9,"Border, Midland and Western"
"Y15-24","IE02",2000,5.5,"Southern and Eastern"
"Y15-24","IS",2000,4.4,"Iceland"
"Y15-24","IS0",2000,4.4,"Ísland"
"Y15-24","IS00",2000,4.4,"Ísland"
"Y15-24","IT",2000,31.5,"Italy"
"Y15-24","ITC",2000,17,"Nord-Ovest"
"Y15-24","ITC1",2000,20.5,"Piemonte"
"Y15-24","ITC2",2000,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",2000,34.9,"Liguria"
"Y15-24","ITC4",2000,13.3,"Lombardia"
"Y15-24","ITF",2000,53.9,"Sud"
"Y15-24","ITF1",2000,26.2,"Abruzzo"
"Y15-24","ITF2",2000,47.2,"Molise"
"Y15-24","ITF3",2000,63.3,"Campania"
"Y15-24","ITF4",2000,45,"Puglia"
"Y15-24","ITF5",2000,40.1,"Basilicata"
"Y15-24","ITF6",2000,64.1,"Calabria"
"Y15-24","ITG",2000,55.8,"Isole"
"Y15-24","ITG1",2000,58,"Sicilia"
"Y15-24","ITG2",2000,49.1,"Sardegna"
"Y15-24","ITH",2000,10.1,"Nord-Est"
"Y15-24","ITH1",2000,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",2000,NA,"Provincia Autonoma di Trento"
"Y15-24","ITH3",2000,9,"Veneto"
"Y15-24","ITH4",2000,8.8,"Friuli-Venezia Giulia"
"Y15-24","ITI",2000,26.9,"Centro (IT)"
"Y15-24","ITI1",2000,17.5,"Toscana"
"Y15-24","ITI2",2000,22.5,"Umbria"
"Y15-24","ITI4",2000,40.2,"Lazio"
"Y15-24","LT",2000,28.6,"Lithuania"
"Y15-24","LT0",2000,28.6,"Lietuva"
"Y15-24","LT00",2000,28.6,"Lietuva"
"Y15-24","LU",2000,6.4,"Luxembourg"
"Y15-24","LU0",2000,6.4,"Luxembourg"
"Y15-24","LU00",2000,6.4,"Luxembourg"
"Y15-24","LV",2000,21.3,"Latvia"
"Y15-24","LV0",2000,21.3,"Latvija"
"Y15-24","LV00",2000,21.3,"Latvija"
"Y15-24","MT",2000,11.8,"Malta"
"Y15-24","MT0",2000,11.8,"Malta"
"Y15-24","MT00",2000,11.8,"Malta"
"Y15-24","NL",2000,5.3,"Netherlands"
"Y15-24","NL1",2000,6.8,"Noord-Nederland"
"Y15-24","NL11",2000,7.3,"Groningen"
"Y15-24","NL12",2000,7.6,"Friesland (NL)"
"Y15-24","NL13",2000,5,"Drenthe"
"Y15-24","NL2",2000,5.1,"Oost-Nederland"
"Y15-24","NL21",2000,5.7,"Overijssel"
"Y15-24","NL22",2000,5.1,"Gelderland"
"Y15-24","NL23",2000,NA,"Flevoland"
"Y15-24","NL3",2000,5.5,"West-Nederland"
"Y15-24","NL31",2000,6.2,"Utrecht"
"Y15-24","NL32",2000,4.2,"Noord-Holland"
"Y15-24","NL33",2000,6.2,"Zuid-Holland"
"Y15-24","NL34",2000,6.1,"Zeeland"
"Y15-24","NL4",2000,4.1,"Zuid-Nederland"
"Y15-24","NL41",2000,3.5,"Noord-Brabant"
"Y15-24","NL42",2000,5.5,"Limburg (NL)"
"Y15-24","NO",2000,11.1,"Norway"
"Y15-24","NO0",2000,11.1,"Norge"
"Y15-24","NO01",2000,8,"Oslo og Akershus"
"Y15-24","NO02",2000,7.2,"Hedmark og Oppland"
"Y15-24","NO03",2000,11.7,"Sør-Østlandet"
"Y15-24","NO04",2000,10.1,"Agder og Rogaland"
"Y15-24","NO05",2000,10.7,"Vestlandet"
"Y15-24","NO06",2000,16.1,"Trøndelag"
"Y15-24","NO07",2000,17.4,"Nord-Norge"
"Y15-24","PL",2000,35.7,"Poland"
"Y15-24","PL1",2000,35.3,"Region Centralny"
"Y15-24","PL11",2000,41.2,"Lódzkie"
"Y15-24","PL12",2000,32,"Mazowieckie"
"Y15-24","PL2",2000,31,"Region Poludniowy"
"Y15-24","PL21",2000,27.6,"Malopolskie"
"Y15-24","PL22",2000,34.1,"Slaskie"
"Y15-24","PL3",2000,37.2,"Region Wschodni"
"Y15-24","PL31",2000,34.9,"Lubelskie"
"Y15-24","PL32",2000,41.6,"Podkarpackie"
"Y15-24","PL33",2000,40.3,"Swietokrzyskie"
"Y15-24","PL34",2000,30.9,"Podlaskie"
"Y15-24","PL4",2000,36.1,"Region Pólnocno-Zachodni"
"Y15-24","PL41",2000,32.9,"Wielkopolskie"
"Y15-24","PL42",2000,46.2,"Zachodniopomorskie"
"Y15-24","PL43",2000,35.4,"Lubuskie"
"Y15-24","PL5",2000,39.3,"Region Poludniowo-Zachodni"
"Y15-24","PL51",2000,42.1,"Dolnoslaskie"
"Y15-24","PL52",2000,31.4,"Opolskie"
"Y15-24","PL6",2000,37.7,"Region Pólnocny"
"Y15-24","PL61",2000,38.1,"Kujawsko-Pomorskie"
"Y15-24","PL62",2000,41.2,"Warminsko-Mazurskie"
"Y15-24","PL63",2000,33.6,"Pomorskie"
"Y15-24","PT",2000,8.2,"Portugal"
"Y15-24","PT1",2000,8.3,"Continente"
"Y15-24","PT11",2000,7.2,"Norte"
"Y15-24","PT15",2000,NA,"Algarve"
"Y15-24","PT16",2000,7.3,"Centro (PT)"
"Y15-24","PT17",2000,10.6,"Área Metropolitana de Lisboa"
"Y15-24","PT18",2000,NA,"Alentejo"
"Y15-24","PT2",2000,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",2000,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",2000,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",2000,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",2000,17.8,"Romania"
"Y15-24","RO1",2000,15.9,"Macroregiunea unu"
"Y15-24","RO11",2000,15.4,"Nord-Vest"
"Y15-24","RO12",2000,16.6,"Centru"
"Y15-24","RO2",2000,17.1,"Macroregiunea doi"
"Y15-24","RO21",2000,15.3,"Nord-Est"
"Y15-24","RO22",2000,20.1,"Sud-Est"
"Y15-24","RO3",2000,21.7,"Macroregiunea trei"
"Y15-24","RO31",2000,21.4,"Sud - Muntenia"
"Y15-24","RO32",2000,22.4,"Bucuresti - Ilfov"
"Y15-24","RO4",2000,17.2,"Macroregiunea patru"
"Y15-24","RO41",2000,14,"Sud-Vest Oltenia"
"Y15-24","RO42",2000,20.9,"Vest"
"Y15-24","SE",2000,9.5,"Sweden"
"Y15-24","SE1",2000,8.5,"Östra Sverige"
"Y15-24","SE11",2000,NA,"Stockholm"
"Y15-24","SE12",2000,NA,"Östra Mellansverige"
"Y15-24","SE2",2000,9.1,"Södra Sverige"
"Y15-24","SE21",2000,NA,"Småland med öarna"
"Y15-24","SE22",2000,15.4,"Sydsverige"
"Y15-24","SE23",2000,NA,"Västsverige"
"Y15-24","SE3",2000,NA,"Norra Sverige"
"Y15-24","SE31",2000,NA,"Norra Mellansverige"
"Y15-24","SE32",2000,NA,"Mellersta Norrland"
"Y15-24","SE33",2000,NA,"Övre Norrland"
"Y15-24","SI",2000,16.4,"Slovenia"
"Y15-24","SI0",2000,16.4,"Slovenija"
"Y15-24","SK",2000,36.9,"Slovakia"
"Y15-24","SK0",2000,36.9,"Slovensko"
"Y15-24","SK01",2000,18.9,"Bratislavský kraj"
"Y15-24","SK02",2000,32.8,"Západné Slovensko"
"Y15-24","SK03",2000,37.5,"Stredné Slovensko"
"Y15-24","SK04",2000,47.4,"Východné Slovensko"
"Y15-24","UK",2000,12,"United Kingdom"
"Y15-24","UKC",2000,20.6,"North East (UK)"
"Y15-24","UKC1",2000,22.1,"Tees Valley and Durham"
"Y15-24","UKC2",2000,19.3,"Northumberland and Tyne and Wear"
"Y15-24","UKD",2000,9.8,"North West (UK)"
"Y15-24","UKD1",2000,NA,"Cumbria"
"Y15-24","UKD3",2000,10.1,"Greater Manchester"
"Y15-24","UKD4",2000,NA,"Lancashire"
"Y15-24","UKE",2000,13.2,"Yorkshire and The Humber"
"Y15-24","UKE1",2000,NA,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",2000,NA,"North Yorkshire"
"Y15-24","UKE3",2000,15.7,"South Yorkshire"
"Y15-24","UKE4",2000,11.2,"West Yorkshire"
"Y15-24","UKF",2000,12.9,"East Midlands (UK)"
"Y15-24","UKF1",2000,13.9,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",2000,11.7,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",2000,NA,"Lincolnshire"
"Y15-24","UKG",2000,13.7,"West Midlands (UK)"
"Y15-24","UKG1",2000,NA,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",2000,10,"Shropshire and Staffordshire"
"Y15-24","UKG3",2000,18.1,"West Midlands"
"Y15-24","UKH",2000,8.7,"East of England"
"Y15-24","UKH1",2000,8.7,"East Anglia"
"Y15-24","UKH2",2000,9,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",2000,NA,"Essex"
"Y15-24","UKI",2000,15.4,"London"
"Y15-24","UKI1",2000,18.4,"Inner London (NUTS 2010)"
"Y15-24","UKI2",2000,13.3,"Outer London (NUTS 2010)"
"Y15-24","UKJ",2000,7.1,"South East (UK)"
"Y15-24","UKJ1",2000,NA,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",2000,6,"Surrey, East and West Sussex"
"Y15-24","UKJ3",2000,8.6,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",2000,10,"Kent"
"Y15-24","UKK",2000,8.9,"South West (UK)"
"Y15-24","UKK1",2000,7.9,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",2000,NA,"Dorset and Somerset"
"Y15-24","UKK3",2000,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",2000,NA,"Devon"
"Y15-24","UKL",2000,14.1,"Wales"
"Y15-24","UKL1",2000,15.1,"West Wales and The Valleys"
"Y15-24","UKL2",2000,NA,"East Wales"
"Y15-24","UKM",2000,15.5,"Scotland"
"Y15-24","UKM2",2000,15,"Eastern Scotland"
"Y15-24","UKM3",2000,18,"South Western Scotland"
"Y15-24","UKM5",2000,NA,"North Eastern Scotland"
"Y15-24","UKM6",2000,NA,"Highlands and Islands"
"Y15-24","UKN",2000,11.4,"Northern Ireland (UK)"
"Y15-24","UKN0",2000,11.4,"Northern Ireland (UK)"
"Y20-64","AT",2000,4.6,"Austria"
"Y20-64","AT1",2000,5.8,"Ostösterreich"
"Y20-64","AT11",2000,4.9,"Burgenland (AT)"
"Y20-64","AT12",2000,4,"Niederösterreich"
"Y20-64","AT13",2000,7.4,"Wien"
"Y20-64","AT2",2000,4.4,"Südösterreich"
"Y20-64","AT21",2000,4.3,"Kärnten"
"Y20-64","AT22",2000,4.5,"Steiermark"
"Y20-64","AT3",2000,3.3,"Westösterreich"
"Y20-64","AT31",2000,3.8,"Oberösterreich"
"Y20-64","AT32",2000,3.2,"Salzburg"
"Y20-64","AT33",2000,2.9,"Tirol"
"Y20-64","AT34",2000,2.7,"Vorarlberg"
"Y20-64","BE",2000,6.3,"Belgium"
"Y20-64","BE1",2000,14.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",2000,14.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",2000,3.4,"Vlaams Gewest"
"Y20-64","BE21",2000,4,"Prov. Antwerpen"
"Y20-64","BE22",2000,4.7,"Prov. Limburg (BE)"
"Y20-64","BE23",2000,3,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",2000,2.7,"Prov. Vlaams-Brabant"
"Y20-64","BE25",2000,2.8,"Prov. West-Vlaanderen"
"Y20-64","BE3",2000,9.6,"Région wallonne"
"Y20-64","BE31",2000,6.7,"Prov. Brabant Wallon"
"Y20-64","BE32",2000,12.1,"Prov. Hainaut"
"Y20-64","BE33",2000,8.1,"Prov. Liège"
"Y20-64","BE34",2000,5.4,"Prov. Luxembourg (BE)"
"Y20-64","BE35",2000,10.7,"Prov. Namur"
"Y20-64","BG",2000,15.8,"Bulgaria"
"Y20-64","BG41",2000,10.8,"Yugozapaden"
"Y20-64","CH",2000,2.5,"Switzerland"
"Y20-64","CH0",2000,2.5,"Schweiz/Suisse/Svizzera"
"Y20-64","CY",2000,4.7,"Cyprus"
"Y20-64","CY0",2000,4.7,"Kypros"
"Y20-64","CY00",2000,4.7,"Kypros"
"Y20-64","CZ",2000,8.4,"Czech Republic"
"Y20-64","CZ0",2000,8.4,"Ceská republika"
"Y20-64","CZ01",2000,3.8,"Praha"
"Y20-64","CZ02",2000,7.4,"Strední Cechy"
"Y20-64","CZ03",2000,5.8,"Jihozápad"
"Y20-64","CZ04",2000,14.2,"Severozápad"
"Y20-64","CZ05",2000,6.6,"Severovýchod"
"Y20-64","CZ06",2000,6.8,"Jihovýchod"
"Y20-64","CZ07",2000,10.4,"Strední Morava"
"Y20-64","CZ08",2000,13.6,"Moravskoslezsko"
"Y20-64","DE",2000,8,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",2000,4.1,"Baden-Württemberg"
"Y20-64","DE11",2000,3.9,"Stuttgart"
"Y20-64","DE12",2000,4.7,"Karlsruhe"
"Y20-64","DE13",2000,4.3,"Freiburg"
"Y20-64","DE14",2000,3.5,"Tübingen"
"Y20-64","DE2",2000,3.9,"Bayern"
"Y20-64","DE21",2000,3,"Oberbayern"
"Y20-64","DE22",2000,3.4,"Niederbayern"
"Y20-64","DE23",2000,4.7,"Oberpfalz"
"Y20-64","DE24",2000,4.8,"Oberfranken"
"Y20-64","DE25",2000,5.7,"Mittelfranken"
"Y20-64","DE26",2000,4.3,"Unterfranken"
"Y20-64","DE27",2000,3.7,"Schwaben"
"Y20-64","DE3",2000,14.4,"Berlin"
"Y20-64","DE30",2000,14.4,"Berlin"
"Y20-64","DE4",2000,16.5,"Brandenburg"
"Y20-64","DE40",2000,16.5,"Brandenburg"
"Y20-64","DE5",2000,10,"Bremen"
"Y20-64","DE50",2000,10,"Bremen"
"Y20-64","DE6",2000,7.8,"Hamburg"
"Y20-64","DE60",2000,7.8,"Hamburg"
"Y20-64","DE7",2000,5.7,"Hessen"
"Y20-64","DE71",2000,5.1,"Darmstadt"
"Y20-64","DE72",2000,6.7,"Gießen"
"Y20-64","DE73",2000,6.9,"Kassel"
"Y20-64","DE8",2000,17,"Mecklenburg-Vorpommern"
"Y20-64","DE80",2000,17,"Mecklenburg-Vorpommern"
"Y20-64","DE9",2000,6.5,"Niedersachsen"
"Y20-64","DE91",2000,7.2,"Braunschweig"
"Y20-64","DE92",2000,7.4,"Hannover"
"Y20-64","DE93",2000,6.2,"Lüneburg"
"Y20-64","DE94",2000,5.5,"Weser-Ems"
"Y20-64","DEA",2000,6.5,"Nordrhein-Westfalen"
"Y20-64","DEA1",2000,6.7,"Düsseldorf"
"Y20-64","DEA2",2000,6.1,"Köln"
"Y20-64","DEA3",2000,5.3,"Münster"
"Y20-64","DEA4",2000,5.6,"Detmold"
"Y20-64","DEA5",2000,7.8,"Arnsberg"
"Y20-64","DEB",2000,5.7,"Rheinland-Pfalz"
"Y20-64","DEC",2000,7.2,"Saarland"
"Y20-64","DEC0",2000,7.2,"Saarland"
"Y20-64","DED",2000,16.5,"Sachsen"
"Y20-64","DED2",2000,16.3,"Dresden"
"Y20-64","DEE",2000,20.8,"Sachsen-Anhalt"
"Y20-64","DEE0",2000,20.8,"Sachsen-Anhalt"
"Y20-64","DEF",2000,6.4,"Schleswig-Holstein"
"Y20-64","DEF0",2000,6.4,"Schleswig-Holstein"
"Y20-64","DEG",2000,13.9,"Thüringen"
"Y20-64","DEG0",2000,13.9,"Thüringen"
"Y20-64","DK",2000,4.3,"Denmark"
"Y20-64","DK0",2000,4.3,"Danmark"
"Y20-64","EA17",2000,9,"Euro area (17 countries)"
"Y20-64","EA18",2000,9.1,"Euro area (18 countries)"
"Y20-64","EA19",2000,9.2,"Euro area (19 countries)"
"Y20-64","EE",2000,13,"Estonia"
"Y20-64","EE0",2000,13,"Eesti"
"Y20-64","EE00",2000,13,"Eesti"
"Y20-64","EL",2000,10.8,"Greece"
"Y20-64","EL1",2000,11,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",2000,8.6,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",2000,10.6,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",2000,14.5,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",2000,12.7,"Thessalia (NUTS 2010)"
"Y20-64","EL2",2000,10.3,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",2000,11.1,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",2000,6,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",2000,10.1,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",2000,13.1,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",2000,9,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",2000,11.8,"Attiki"
"Y20-64","EL30",2000,11.8,"Attiki"
"Y20-64","EL4",2000,7.8,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",2000,7.7,"Voreio Aigaio"
"Y20-64","EL42",2000,10.1,"Notio Aigaio"
"Y20-64","EL43",2000,6.8,"Kriti"
"Y20-64","ES",2000,13.2,"Spain"
"Y20-64","ES1",2000,14.9,"Noroeste (ES)"
"Y20-64","ES11",2000,14.4,"Galicia"
"Y20-64","ES12",2000,17.1,"Principado de Asturias"
"Y20-64","ES13",2000,13.2,"Cantabria"
"Y20-64","ES2",2000,9,"Noreste (ES)"
"Y20-64","ES21",2000,11.7,"País Vasco"
"Y20-64","ES22",2000,4.1,"Comunidad Foral de Navarra"
"Y20-64","ES23",2000,7.7,"La Rioja"
"Y20-64","ES24",2000,6.7,"Aragón"
"Y20-64","ES3",2000,11.1,"Comunidad de Madrid"
"Y20-64","ES30",2000,11.1,"Comunidad de Madrid"
"Y20-64","ES4",2000,14.8,"Centro (ES)"
"Y20-64","ES41",2000,13.1,"Castilla y León"
"Y20-64","ES42",2000,11.7,"Castilla-la Mancha"
"Y20-64","ES43",2000,23.4,"Extremadura"
"Y20-64","ES5",2000,8.7,"Este (ES)"
"Y20-64","ES51",2000,8,"Cataluña"
"Y20-64","ES52",2000,10.8,"Comunidad Valenciana"
"Y20-64","ES53",2000,4.6,"Illes Balears"
"Y20-64","ES6",2000,21.6,"Sur (ES)"
"Y20-64","ES61",2000,23.4,"Andalucía"
"Y20-64","ES62",2000,10.7,"Región de Murcia"
"Y20-64","ES63",2000,24.4,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",2000,20.9,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",2000,13.4,"Canarias (ES)"
"Y20-64","ES70",2000,13.4,"Canarias (ES)"
"Y20-64","EU15",2000,8.1,"European Union (15 countries)"
"Y20-64","EU27",2000,9,"European Union (27 countries)"
"Y20-64","FI",2000,9.2,"Finland"
"Y20-64","FI1",2000,9.2,"Manner-Suomi"
"Y20-64","FI19",2000,9.6,"Länsi-Suomi"
"Y20-64","FI2",2000,NA,"Åland"
"Y20-64","FI20",2000,NA,"Åland"
"Y20-64","FR",2000,9.9,"France"
"Y20-64","FR1",2000,8.5,"Île de France"
"Y20-64","FR10",2000,8.5,"Île de France"
"Y20-64","FR2",2000,9.6,"Bassin Parisien"
"Y20-64","FR21",2000,10.9,"Champagne-Ardenne"
"Y20-64","FR22",2000,11,"Picardie"
"Y20-64","FR23",2000,10.6,"Haute-Normandie"
"Y20-64","FR24",2000,8.1,"Centre (FR)"
"Y20-64","FR25",2000,8.1,"Basse-Normandie"
"Y20-64","FR26",2000,9.2,"Bourgogne"
"Y20-64","FR3",2000,15.9,"Nord - Pas-de-Calais"
"Y20-64","FR30",2000,15.9,"Nord - Pas-de-Calais"
"Y20-64","FR4",2000,8,"Est (FR)"
"Y20-64","FR41",2000,9.5,"Lorraine"
"Y20-64","FR42",2000,6.3,"Alsace"
"Y20-64","FR43",2000,7.6,"Franche-Comté"
"Y20-64","FR5",2000,8.3,"Ouest (FR)"
"Y20-64","FR51",2000,9.3,"Pays de la Loire"
"Y20-64","FR52",2000,7.2,"Bretagne"
"Y20-64","FR53",2000,8.2,"Poitou-Charentes"
"Y20-64","FR6",2000,10,"Sud-Ouest (FR)"
"Y20-64","FR61",2000,10.7,"Aquitaine"
"Y20-64","FR62",2000,9.7,"Midi-Pyrénées"
"Y20-64","FR63",2000,7.5,"Limousin"
"Y20-64","FR7",2000,8.3,"Centre-Est (FR)"
"Y20-64","FR71",2000,8,"Rhône-Alpes"
"Y20-64","FR72",2000,9.9,"Auvergne"
"Y20-64","FR8",2000,15,"Méditerranée"
"Y20-64","FR81",2000,16.2,"Languedoc-Roussillon"
"Y20-64","FR82",2000,14.1,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",2000,21.8,"Corse"
"Y20-64","HU",2000,6.3,"Hungary"
"Y20-64","HU1",2000,5.3,"Közép-Magyarország"
"Y20-64","HU10",2000,5.3,"Közép-Magyarország"
"Y20-64","HU2",2000,5.5,"Dunántúl"
"Y20-64","HU21",2000,5,"Közép-Dunántúl"
"Y20-64","HU22",2000,4.2,"Nyugat-Dunántúl"
"Y20-64","HU23",2000,7.7,"Dél-Dunántúl"
"Y20-64","HU3",2000,7.8,"Alföld és Észak"
"Y20-64","HU31",2000,9.6,"Észak-Magyarország"
"Y20-64","HU32",2000,9.3,"Észak-Alföld"
"Y20-64","HU33",2000,4.7,"Dél-Alföld"
"Y20-64","IE",2000,4,"Ireland"
"Y20-64","IE0",2000,4,"Éire/Ireland"
"Y20-64","IE01",2000,5.3,"Border, Midland and Western"
"Y20-64","IE02",2000,3.6,"Southern and Eastern"
"Y20-64","IS",2000,1.5,"Iceland"
"Y20-64","IS0",2000,1.5,"Ísland"
"Y20-64","IS00",2000,1.5,"Ísland"
"Y20-64","IT",2000,10.3,"Italy"
"Y20-64","ITC",2000,5.1,"Nord-Ovest"
"Y20-64","ITC1",2000,6.1,"Piemonte"
"Y20-64","ITC2",2000,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",2000,8.8,"Liguria"
"Y20-64","ITC4",2000,4,"Lombardia"
"Y20-64","ITF",2000,19.2,"Sud"
"Y20-64","ITF1",2000,7.3,"Abruzzo"
"Y20-64","ITF2",2000,12.8,"Molise"
"Y20-64","ITF3",2000,22.2,"Campania"
"Y20-64","ITF4",2000,16.4,"Puglia"
"Y20-64","ITF5",2000,16.4,"Basilicata"
"Y20-64","ITF6",2000,26.1,"Calabria"
"Y20-64","ITG",2000,22,"Isole"
"Y20-64","ITG1",2000,22.9,"Sicilia"
"Y20-64","ITG2",2000,19.4,"Sardegna"
"Y20-64","ITH",2000,4,"Nord-Est"
"Y20-64","ITH1",2000,2.3,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",2000,3.2,"Provincia Autonoma di Trento"
"Y20-64","ITH3",2000,3.9,"Veneto"
"Y20-64","ITH4",2000,4,"Friuli-Venezia Giulia"
"Y20-64","ITI",2000,8.6,"Centro (IT)"
"Y20-64","ITI1",2000,6.5,"Toscana"
"Y20-64","ITI2",2000,6.3,"Umbria"
"Y20-64","ITI4",2000,11.3,"Lazio"
"Y20-64","LT",2000,15.9,"Lithuania"
"Y20-64","LT0",2000,15.9,"Lietuva"
"Y20-64","LT00",2000,15.9,"Lietuva"
"Y20-64","LU",2000,2.3,"Luxembourg"
"Y20-64","LU0",2000,2.3,"Luxembourg"
"Y20-64","LU00",2000,2.3,"Luxembourg"
"Y20-64","LV",2000,14,"Latvia"
"Y20-64","LV0",2000,14,"Latvija"
"Y20-64","LV00",2000,14,"Latvija"
"Y20-64","MT",2000,4.8,"Malta"
"Y20-64","MT0",2000,4.8,"Malta"
"Y20-64","MT00",2000,4.8,"Malta"
"Y20-64","NL",2000,2.3,"Netherlands"
"Y20-64","NL1",2000,3.5,"Noord-Nederland"
"Y20-64","NL11",2000,3.7,"Groningen"
"Y20-64","NL12",2000,3.7,"Friesland (NL)"
"Y20-64","NL13",2000,3,"Drenthe"
"Y20-64","NL2",2000,2.2,"Oost-Nederland"
"Y20-64","NL21",2000,2.2,"Overijssel"
"Y20-64","NL22",2000,2,"Gelderland"
"Y20-64","NL23",2000,3.6,"Flevoland"
"Y20-64","NL3",2000,2.3,"West-Nederland"
"Y20-64","NL31",2000,1.8,"Utrecht"
"Y20-64","NL32",2000,2.6,"Noord-Holland"
"Y20-64","NL33",2000,2.3,"Zuid-Holland"
"Y20-64","NL34",2000,2.7,"Zeeland"
"Y20-64","NL4",2000,2,"Zuid-Nederland"
"Y20-64","NL41",2000,1.8,"Noord-Brabant"
"Y20-64","NL42",2000,2.3,"Limburg (NL)"
"Y20-64","NO",2000,2.6,"Norway"
"Y20-64","NO0",2000,2.6,"Norge"
"Y20-64","NO01",2000,1.9,"Oslo og Akershus"
"Y20-64","NO02",2000,2.3,"Hedmark og Oppland"
"Y20-64","NO03",2000,2.5,"Sør-Østlandet"
"Y20-64","NO04",2000,3.6,"Agder og Rogaland"
"Y20-64","NO05",2000,2.7,"Vestlandet"
"Y20-64","NO06",2000,3.1,"Trøndelag"
"Y20-64","NO07",2000,3,"Nord-Norge"
"Y20-64","PL",2000,16.3,"Poland"
"Y20-64","PL1",2000,14.4,"Region Centralny"
"Y20-64","PL11",2000,16.1,"Lódzkie"
"Y20-64","PL12",2000,13.3,"Mazowieckie"
"Y20-64","PL2",2000,15.2,"Region Poludniowy"
"Y20-64","PL21",2000,11.8,"Malopolskie"
"Y20-64","PL22",2000,18.4,"Slaskie"
"Y20-64","PL3",2000,15.1,"Region Wschodni"
"Y20-64","PL31",2000,14,"Lubelskie"
"Y20-64","PL32",2000,14.7,"Podkarpackie"
"Y20-64","PL33",2000,17.3,"Swietokrzyskie"
"Y20-64","PL34",2000,15.9,"Podlaskie"
"Y20-64","PL4",2000,16.5,"Region Pólnocno-Zachodni"
"Y20-64","PL41",2000,13.9,"Wielkopolskie"
"Y20-64","PL42",2000,19.8,"Zachodniopomorskie"
"Y20-64","PL43",2000,21,"Lubuskie"
"Y20-64","PL5",2000,20.4,"Region Poludniowo-Zachodni"
"Y20-64","PL51",2000,22.6,"Dolnoslaskie"
"Y20-64","PL52",2000,14.7,"Opolskie"
"Y20-64","PL6",2000,18.7,"Region Pólnocny"
"Y20-64","PL61",2000,18,"Kujawsko-Pomorskie"
"Y20-64","PL62",2000,21.8,"Warminsko-Mazurskie"
"Y20-64","PL63",2000,16.8,"Pomorskie"
"Y20-64","PT",2000,3.8,"Portugal"
"Y20-64","PT1",2000,3.9,"Continente"
"Y20-64","PT11",2000,3.9,"Norte"
"Y20-64","PT15",2000,NA,"Algarve"
"Y20-64","PT16",2000,1.9,"Centro (PT)"
"Y20-64","PT17",2000,5.2,"Área Metropolitana de Lisboa"
"Y20-64","PT18",2000,5.5,"Alentejo"
"Y20-64","PT2",2000,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",2000,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",2000,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",2000,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",2000,7.1,"Romania"
"Y20-64","RO1",2000,7.2,"Macroregiunea unu"
"Y20-64","RO11",2000,7.1,"Nord-Vest"
"Y20-64","RO12",2000,7.4,"Centru"
"Y20-64","RO2",2000,8.1,"Macroregiunea doi"
"Y20-64","RO21",2000,7.4,"Nord-Est"
"Y20-64","RO22",2000,9,"Sud-Est"
"Y20-64","RO3",2000,6.6,"Macroregiunea trei"
"Y20-64","RO31",2000,6.7,"Sud - Muntenia"
"Y20-64","RO32",2000,6.5,"Bucuresti - Ilfov"
"Y20-64","RO4",2000,6.2,"Macroregiunea patru"
"Y20-64","RO41",2000,5.3,"Sud-Vest Oltenia"
"Y20-64","RO42",2000,7.4,"Vest"
"Y20-64","SE",2000,5.4,"Sweden"
"Y20-64","SE1",2000,4.1,"Östra Sverige"
"Y20-64","SE11",2000,3.2,"Stockholm"
"Y20-64","SE12",2000,5.4,"Östra Mellansverige"
"Y20-64","SE2",2000,5.6,"Södra Sverige"
"Y20-64","SE21",2000,4.4,"Småland med öarna"
"Y20-64","SE22",2000,7,"Sydsverige"
"Y20-64","SE23",2000,5.2,"Västsverige"
"Y20-64","SE3",2000,7.7,"Norra Sverige"
"Y20-64","SE31",2000,6.7,"Norra Mellansverige"
"Y20-64","SE32",2000,8,"Mellersta Norrland"
"Y20-64","SE33",2000,9.1,"Övre Norrland"
"Y20-64","SI",2000,6.7,"Slovenia"
"Y20-64","SI0",2000,6.7,"Slovenija"
"Y20-64","SK",2000,17.6,"Slovakia"
"Y20-64","SK0",2000,17.6,"Slovensko"
"Y20-64","SK01",2000,6.6,"Bratislavský kraj"
"Y20-64","SK02",2000,16.5,"Západné Slovensko"
"Y20-64","SK03",2000,19.5,"Stredné Slovensko"
"Y20-64","SK04",2000,22.7,"Východné Slovensko"
"Y20-64","UK",2000,5,"United Kingdom"
"Y20-64","UKC",2000,7.8,"North East (UK)"
"Y20-64","UKC1",2000,7.6,"Tees Valley and Durham"
"Y20-64","UKC2",2000,8,"Northumberland and Tyne and Wear"
"Y20-64","UKD",2000,4.9,"North West (UK)"
"Y20-64","UKD1",2000,NA,"Cumbria"
"Y20-64","UKD3",2000,4.5,"Greater Manchester"
"Y20-64","UKD4",2000,4.1,"Lancashire"
"Y20-64","UKE",2000,5,"Yorkshire and The Humber"
"Y20-64","UKE1",2000,6,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",2000,3.7,"North Yorkshire"
"Y20-64","UKE3",2000,5.8,"South Yorkshire"
"Y20-64","UKE4",2000,4.7,"West Yorkshire"
"Y20-64","UKF",2000,4.4,"East Midlands (UK)"
"Y20-64","UKF1",2000,5,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",2000,4.1,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",2000,3.6,"Lincolnshire"
"Y20-64","UKG",2000,5.3,"West Midlands (UK)"
"Y20-64","UKG1",2000,3.8,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",2000,3.9,"Shropshire and Staffordshire"
"Y20-64","UKG3",2000,7,"West Midlands"
"Y20-64","UKH",2000,3.1,"East of England"
"Y20-64","UKH1",2000,3.8,"East Anglia"
"Y20-64","UKH2",2000,2.4,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",2000,3,"Essex"
"Y20-64","UKI",2000,6.5,"London"
"Y20-64","UKI1",2000,8.7,"Inner London (NUTS 2010)"
"Y20-64","UKI2",2000,5.1,"Outer London (NUTS 2010)"
"Y20-64","UKJ",2000,3.2,"South East (UK)"
"Y20-64","UKJ1",2000,2,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",2000,3,"Surrey, East and West Sussex"
"Y20-64","UKJ3",2000,3.7,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",2000,4.8,"Kent"
"Y20-64","UKK",2000,3.7,"South West (UK)"
"Y20-64","UKK1",2000,2.6,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",2000,4.3,"Dorset and Somerset"
"Y20-64","UKK3",2000,6.4,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",2000,4.5,"Devon"
"Y20-64","UKL",2000,5.6,"Wales"
"Y20-64","UKL1",2000,6.1,"West Wales and The Valleys"
"Y20-64","UKL2",2000,4.8,"East Wales"
"Y20-64","UKM",2000,6.7,"Scotland"
"Y20-64","UKM2",2000,5.9,"Eastern Scotland"
"Y20-64","UKM3",2000,8.3,"South Western Scotland"
"Y20-64","UKM5",2000,NA,"North Eastern Scotland"
"Y20-64","UKM6",2000,7.2,"Highlands and Islands"
"Y20-64","UKN",2000,6.6,"Northern Ireland (UK)"
"Y20-64","UKN0",2000,6.6,"Northern Ireland (UK)"
"Y_GE15","AT",2000,4.7,"Austria"
"Y_GE15","AT1",2000,5.8,"Ostösterreich"
"Y_GE15","AT11",2000,4.8,"Burgenland (AT)"
"Y_GE15","AT12",2000,4.1,"Niederösterreich"
"Y_GE15","AT13",2000,7.5,"Wien"
"Y_GE15","AT2",2000,4.6,"Südösterreich"
"Y_GE15","AT21",2000,4.6,"Kärnten"
"Y_GE15","AT22",2000,4.5,"Steiermark"
"Y_GE15","AT3",2000,3.5,"Westösterreich"
"Y_GE15","AT31",2000,3.9,"Oberösterreich"
"Y_GE15","AT32",2000,3.3,"Salzburg"
"Y_GE15","AT33",2000,3,"Tirol"
"Y_GE15","AT34",2000,2.8,"Vorarlberg"
"Y_GE15","BE",2000,6.6,"Belgium"
"Y_GE15","BE1",2000,14.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",2000,14.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",2000,3.6,"Vlaams Gewest"
"Y_GE15","BE21",2000,4.3,"Prov. Antwerpen"
"Y_GE15","BE22",2000,5.1,"Prov. Limburg (BE)"
"Y_GE15","BE23",2000,3.1,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",2000,2.9,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",2000,3,"Prov. West-Vlaanderen"
"Y_GE15","BE3",2000,9.8,"Région wallonne"
"Y_GE15","BE31",2000,7.2,"Prov. Brabant Wallon"
"Y_GE15","BE32",2000,12.3,"Prov. Hainaut"
"Y_GE15","BE33",2000,8.4,"Prov. Liège"
"Y_GE15","BE34",2000,5.5,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",2000,10.8,"Prov. Namur"
"Y_GE15","BG",2000,16.2,"Bulgaria"
"Y_GE15","BG41",2000,11.1,"Yugozapaden"
"Y_GE15","CH",2000,2.7,"Switzerland"
"Y_GE15","CH0",2000,2.7,"Schweiz/Suisse/Svizzera"
"Y_GE15","CY",2000,5,"Cyprus"
"Y_GE15","CY0",2000,5,"Kypros"
"Y_GE15","CY00",2000,5,"Kypros"
"Y_GE15","CZ",2000,8.8,"Czech Republic"
"Y_GE15","CZ0",2000,8.8,"Ceská republika"
"Y_GE15","CZ01",2000,4,"Praha"
"Y_GE15","CZ02",2000,7.5,"Strední Cechy"
"Y_GE15","CZ03",2000,6,"Jihozápad"
"Y_GE15","CZ04",2000,15,"Severozápad"
"Y_GE15","CZ05",2000,6.8,"Severovýchod"
"Y_GE15","CZ06",2000,7.1,"Jihovýchod"
"Y_GE15","CZ07",2000,10.9,"Strední Morava"
"Y_GE15","CZ08",2000,14.1,"Moravskoslezsko"
"Y_GE15","DE",2000,7.9,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",2000,4.1,"Baden-Württemberg"
"Y_GE15","DE11",2000,3.9,"Stuttgart"
"Y_GE15","DE12",2000,4.7,"Karlsruhe"
"Y_GE15","DE13",2000,4.4,"Freiburg"
"Y_GE15","DE14",2000,3.5,"Tübingen"
"Y_GE15","DE2",2000,4,"Bayern"
"Y_GE15","DE21",2000,3,"Oberbayern"
"Y_GE15","DE22",2000,3.3,"Niederbayern"
"Y_GE15","DE23",2000,4.6,"Oberpfalz"
"Y_GE15","DE24",2000,4.9,"Oberfranken"
"Y_GE15","DE25",2000,5.6,"Mittelfranken"
"Y_GE15","DE26",2000,4.5,"Unterfranken"
"Y_GE15","DE27",2000,3.8,"Schwaben"
"Y_GE15","DE3",2000,14.4,"Berlin"
"Y_GE15","DE30",2000,14.4,"Berlin"
"Y_GE15","DE4",2000,16.3,"Brandenburg"
"Y_GE15","DE40",2000,16.3,"Brandenburg"
"Y_GE15","DE5",2000,10,"Bremen"
"Y_GE15","DE50",2000,10,"Bremen"
"Y_GE15","DE6",2000,7.8,"Hamburg"
"Y_GE15","DE60",2000,7.8,"Hamburg"
"Y_GE15","DE7",2000,5.8,"Hessen"
"Y_GE15","DE71",2000,5.2,"Darmstadt"
"Y_GE15","DE72",2000,6.6,"Gießen"
"Y_GE15","DE73",2000,6.9,"Kassel"
"Y_GE15","DE8",2000,16.4,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",2000,16.4,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",2000,6.6,"Niedersachsen"
"Y_GE15","DE91",2000,7.4,"Braunschweig"
"Y_GE15","DE92",2000,7.4,"Hannover"
"Y_GE15","DE93",2000,6.2,"Lüneburg"
"Y_GE15","DE94",2000,5.5,"Weser-Ems"
"Y_GE15","DEA",2000,6.5,"Nordrhein-Westfalen"
"Y_GE15","DEA1",2000,6.8,"Düsseldorf"
"Y_GE15","DEA2",2000,6,"Köln"
"Y_GE15","DEA3",2000,5.4,"Münster"
"Y_GE15","DEA4",2000,5.7,"Detmold"
"Y_GE15","DEA5",2000,7.7,"Arnsberg"
"Y_GE15","DEB",2000,5.8,"Rheinland-Pfalz"
"Y_GE15","DEC",2000,7.3,"Saarland"
"Y_GE15","DEC0",2000,7.3,"Saarland"
"Y_GE15","DED",2000,16.1,"Sachsen"
"Y_GE15","DED2",2000,15.9,"Dresden"
"Y_GE15","DEE",2000,20.2,"Sachsen-Anhalt"
"Y_GE15","DEE0",2000,20.2,"Sachsen-Anhalt"
"Y_GE15","DEF",2000,6.4,"Schleswig-Holstein"
"Y_GE15","DEF0",2000,6.4,"Schleswig-Holstein"
"Y_GE15","DEG",2000,13.5,"Thüringen"
"Y_GE15","DEG0",2000,13.5,"Thüringen"
"Y_GE15","DK",2000,4.5,"Denmark"
"Y_GE15","DK0",2000,4.5,"Danmark"
"Y_GE15","EA17",2000,9.3,"Euro area (17 countries)"
"Y_GE15","EA18",2000,9.4,"Euro area (18 countries)"
"Y_GE15","EA19",2000,9.4,"Euro area (19 countries)"
"Y_GE15","EE",2000,13.4,"Estonia"
"Y_GE15","EE0",2000,13.4,"Eesti"
"Y_GE15","EE00",2000,13.4,"Eesti"
"Y_GE15","EL",2000,11.2,"Greece"
"Y_GE15","EL1",2000,11.3,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",2000,8.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",2000,10.9,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",2000,15,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",2000,13,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",2000,10.8,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",2000,10.9,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",2000,5.6,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",2000,10.6,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",2000,14.4,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",2000,9.7,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",2000,12.3,"Attiki"
"Y_GE15","EL30",2000,12.3,"Attiki"
"Y_GE15","EL4",2000,8.2,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",2000,7.7,"Voreio Aigaio"
"Y_GE15","EL42",2000,10.5,"Notio Aigaio"
"Y_GE15","EL43",2000,7.2,"Kriti"
"Y_GE15","ES",2000,13.8,"Spain"
"Y_GE15","ES1",2000,15.1,"Noroeste (ES)"
"Y_GE15","ES11",2000,14.7,"Galicia"
"Y_GE15","ES12",2000,17.3,"Principado de Asturias"
"Y_GE15","ES13",2000,13.4,"Cantabria"
"Y_GE15","ES2",2000,9.3,"Noreste (ES)"
"Y_GE15","ES21",2000,11.9,"País Vasco"
"Y_GE15","ES22",2000,4.5,"Comunidad Foral de Navarra"
"Y_GE15","ES23",2000,7.9,"La Rioja"
"Y_GE15","ES24",2000,7,"Aragón"
"Y_GE15","ES3",2000,11.6,"Comunidad de Madrid"
"Y_GE15","ES30",2000,11.6,"Comunidad de Madrid"
"Y_GE15","ES4",2000,15.3,"Centro (ES)"
"Y_GE15","ES41",2000,13.7,"Castilla y León"
"Y_GE15","ES42",2000,12.2,"Castilla-la Mancha"
"Y_GE15","ES43",2000,24.2,"Extremadura"
"Y_GE15","ES5",2000,9.4,"Este (ES)"
"Y_GE15","ES51",2000,8.8,"Cataluña"
"Y_GE15","ES52",2000,11.4,"Comunidad Valenciana"
"Y_GE15","ES53",2000,5.3,"Illes Balears"
"Y_GE15","ES6",2000,22.4,"Sur (ES)"
"Y_GE15","ES61",2000,24.2,"Andalucía"
"Y_GE15","ES62",2000,11.4,"Región de Murcia"
"Y_GE15","ES63",2000,26,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",2000,21.2,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",2000,13.9,"Canarias (ES)"
"Y_GE15","ES70",2000,13.9,"Canarias (ES)"
"Y_GE15","EU15",2000,8.4,"European Union (15 countries)"
"Y_GE15","EU27",2000,9.2,"European Union (27 countries)"
"Y_GE15","FI",2000,11.1,"Finland"
"Y_GE15","FI1",2000,11.2,"Manner-Suomi"
"Y_GE15","FI19",2000,11.5,"Länsi-Suomi"
"Y_GE15","FI2",2000,NA,"Åland"
"Y_GE15","FI20",2000,NA,"Åland"
"Y_GE15","FR",2000,10.2,"France"
"Y_GE15","FR1",2000,8.7,"Île de France"
"Y_GE15","FR10",2000,8.7,"Île de France"
"Y_GE15","FR2",2000,9.9,"Bassin Parisien"
"Y_GE15","FR21",2000,11.3,"Champagne-Ardenne"
"Y_GE15","FR22",2000,11.6,"Picardie"
"Y_GE15","FR23",2000,11,"Haute-Normandie"
"Y_GE15","FR24",2000,8.2,"Centre (FR)"
"Y_GE15","FR25",2000,8.2,"Basse-Normandie"
"Y_GE15","FR26",2000,9.3,"Bourgogne"
"Y_GE15","FR3",2000,16.7,"Nord - Pas-de-Calais"
"Y_GE15","FR30",2000,16.7,"Nord - Pas-de-Calais"
"Y_GE15","FR4",2000,8.3,"Est (FR)"
"Y_GE15","FR41",2000,9.7,"Lorraine"
"Y_GE15","FR42",2000,6.5,"Alsace"
"Y_GE15","FR43",2000,8.1,"Franche-Comté"
"Y_GE15","FR5",2000,8.6,"Ouest (FR)"
"Y_GE15","FR51",2000,9.5,"Pays de la Loire"
"Y_GE15","FR52",2000,7.5,"Bretagne"
"Y_GE15","FR53",2000,8.4,"Poitou-Charentes"
"Y_GE15","FR6",2000,10.3,"Sud-Ouest (FR)"
"Y_GE15","FR61",2000,11.1,"Aquitaine"
"Y_GE15","FR62",2000,10.1,"Midi-Pyrénées"
"Y_GE15","FR63",2000,7.8,"Limousin"
"Y_GE15","FR7",2000,8.5,"Centre-Est (FR)"
"Y_GE15","FR71",2000,8.1,"Rhône-Alpes"
"Y_GE15","FR72",2000,10.2,"Auvergne"
"Y_GE15","FR8",2000,15.3,"Méditerranée"
"Y_GE15","FR81",2000,16.6,"Languedoc-Roussillon"
"Y_GE15","FR82",2000,14.3,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",2000,22.8,"Corse"
"Y_GE15","HU",2000,6.6,"Hungary"
"Y_GE15","HU1",2000,5.5,"Közép-Magyarország"
"Y_GE15","HU10",2000,5.5,"Közép-Magyarország"
"Y_GE15","HU2",2000,5.7,"Dunántúl"
"Y_GE15","HU21",2000,5.2,"Közép-Dunántúl"
"Y_GE15","HU22",2000,4.4,"Nyugat-Dunántúl"
"Y_GE15","HU23",2000,7.9,"Dél-Dunántúl"
"Y_GE15","HU3",2000,8.2,"Alföld és Észak"
"Y_GE15","HU31",2000,10,"Észak-Magyarország"
"Y_GE15","HU32",2000,9.7,"Észak-Alföld"
"Y_GE15","HU33",2000,5,"Dél-Alföld"
"Y_GE15","IE",2000,4.3,"Ireland"
"Y_GE15","IE0",2000,4.3,"Éire/Ireland"
"Y_GE15","IE01",2000,5.7,"Border, Midland and Western"
"Y_GE15","IE02",2000,3.9,"Southern and Eastern"
"Y_GE15","IS",2000,1.9,"Iceland"
"Y_GE15","IS0",2000,1.9,"Ísland"
"Y_GE15","IS00",2000,1.9,"Ísland"
"Y_GE15","IT",2000,10.8,"Italy"
"Y_GE15","ITC",2000,5.5,"Nord-Ovest"
"Y_GE15","ITC1",2000,6.6,"Piemonte"
"Y_GE15","ITC2",2000,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",2000,9.2,"Liguria"
"Y_GE15","ITC4",2000,4.4,"Lombardia"
"Y_GE15","ITF",2000,20.1,"Sud"
"Y_GE15","ITF1",2000,7.5,"Abruzzo"
"Y_GE15","ITF2",2000,13.4,"Molise"
"Y_GE15","ITF3",2000,23.3,"Campania"
"Y_GE15","ITF4",2000,17.3,"Puglia"
"Y_GE15","ITF5",2000,17.1,"Basilicata"
"Y_GE15","ITF6",2000,27.3,"Calabria"
"Y_GE15","ITG",2000,22.9,"Isole"
"Y_GE15","ITG1",2000,23.9,"Sicilia"
"Y_GE15","ITG2",2000,20.2,"Sardegna"
"Y_GE15","ITH",2000,4.2,"Nord-Est"
"Y_GE15","ITH1",2000,2.4,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",2000,3.7,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",2000,4.1,"Veneto"
"Y_GE15","ITH4",2000,4.2,"Friuli-Venezia Giulia"
"Y_GE15","ITI",2000,8.8,"Centro (IT)"
"Y_GE15","ITI1",2000,6.6,"Toscana"
"Y_GE15","ITI2",2000,6.6,"Umbria"
"Y_GE15","ITI4",2000,11.7,"Lazio"
"Y_GE15","LT",2000,15.9,"Lithuania"
"Y_GE15","LT0",2000,15.9,"Lietuva"
"Y_GE15","LT00",2000,15.9,"Lietuva"
"Y_GE15","LU",2000,2.3,"Luxembourg"
"Y_GE15","LU0",2000,2.3,"Luxembourg"
"Y_GE15","LU00",2000,2.3,"Luxembourg"
"Y_GE15","LV",2000,14.2,"Latvia"
"Y_GE15","LV0",2000,14.2,"Latvija"
"Y_GE15","LV00",2000,14.2,"Latvija"
"Y_GE15","MT",2000,6.3,"Malta"
"Y_GE15","MT0",2000,6.3,"Malta"
"Y_GE15","MT00",2000,6.3,"Malta"
"Y_GE15","NL",2000,2.7,"Netherlands"
"Y_GE15","NL1",2000,4.2,"Noord-Nederland"
"Y_GE15","NL11",2000,4.4,"Groningen"
"Y_GE15","NL12",2000,4.5,"Friesland (NL)"
"Y_GE15","NL13",2000,3.5,"Drenthe"
"Y_GE15","NL2",2000,2.7,"Oost-Nederland"
"Y_GE15","NL21",2000,2.6,"Overijssel"
"Y_GE15","NL22",2000,2.5,"Gelderland"
"Y_GE15","NL23",2000,3.8,"Flevoland"
"Y_GE15","NL3",2000,2.6,"West-Nederland"
"Y_GE15","NL31",2000,2.1,"Utrecht"
"Y_GE15","NL32",2000,2.7,"Noord-Holland"
"Y_GE15","NL33",2000,2.7,"Zuid-Holland"
"Y_GE15","NL34",2000,3.4,"Zeeland"
"Y_GE15","NL4",2000,2.3,"Zuid-Nederland"
"Y_GE15","NL41",2000,2.1,"Noord-Brabant"
"Y_GE15","NL42",2000,2.7,"Limburg (NL)"
"Y_GE15","NO",2000,3.5,"Norway"
"Y_GE15","NO0",2000,3.5,"Norge"
"Y_GE15","NO01",2000,2.6,"Oslo og Akershus"
"Y_GE15","NO02",2000,2.7,"Hedmark og Oppland"
"Y_GE15","NO03",2000,3.3,"Sør-Østlandet"
"Y_GE15","NO04",2000,4.1,"Agder og Rogaland"
"Y_GE15","NO05",2000,3.6,"Vestlandet"
"Y_GE15","NO06",2000,4.1,"Trøndelag"
"Y_GE15","NO07",2000,4.5,"Nord-Norge"
"Y_GE15","PL",2000,16.3,"Poland"
"Y_GE15","PL1",2000,14.4,"Region Centralny"
"Y_GE15","PL11",2000,16.2,"Lódzkie"
"Y_GE15","PL12",2000,13.3,"Mazowieckie"
"Y_GE15","PL2",2000,15.4,"Region Poludniowy"
"Y_GE15","PL21",2000,11.6,"Malopolskie"
"Y_GE15","PL22",2000,18.9,"Slaskie"
"Y_GE15","PL3",2000,14.8,"Region Wschodni"
"Y_GE15","PL31",2000,13.6,"Lubelskie"
"Y_GE15","PL32",2000,14.5,"Podkarpackie"
"Y_GE15","PL33",2000,16.9,"Swietokrzyskie"
"Y_GE15","PL34",2000,15.7,"Podlaskie"
"Y_GE15","PL4",2000,16.9,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",2000,14.1,"Wielkopolskie"
"Y_GE15","PL42",2000,20.4,"Zachodniopomorskie"
"Y_GE15","PL43",2000,21.3,"Lubuskie"
"Y_GE15","PL5",2000,20.4,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",2000,22.6,"Dolnoslaskie"
"Y_GE15","PL52",2000,14.6,"Opolskie"
"Y_GE15","PL6",2000,19,"Region Pólnocny"
"Y_GE15","PL61",2000,18.2,"Kujawsko-Pomorskie"
"Y_GE15","PL62",2000,22.4,"Warminsko-Mazurskie"
"Y_GE15","PL63",2000,17.1,"Pomorskie"
"Y_GE15","PT",2000,3.8,"Portugal"
"Y_GE15","PT1",2000,3.9,"Continente"
"Y_GE15","PT11",2000,3.9,"Norte"
"Y_GE15","PT15",2000,NA,"Algarve"
"Y_GE15","PT16",2000,1.9,"Centro (PT)"
"Y_GE15","PT17",2000,5.4,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",2000,5.6,"Alentejo"
"Y_GE15","PT2",2000,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",2000,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",2000,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",2000,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",2000,7,"Romania"
"Y_GE15","RO1",2000,7.2,"Macroregiunea unu"
"Y_GE15","RO11",2000,7,"Nord-Vest"
"Y_GE15","RO12",2000,7.4,"Centru"
"Y_GE15","RO2",2000,7.7,"Macroregiunea doi"
"Y_GE15","RO21",2000,6.8,"Nord-Est"
"Y_GE15","RO22",2000,8.9,"Sud-Est"
"Y_GE15","RO3",2000,6.6,"Macroregiunea trei"
"Y_GE15","RO31",2000,6.6,"Sud - Muntenia"
"Y_GE15","RO32",2000,6.6,"Bucuresti - Ilfov"
"Y_GE15","RO4",2000,6.1,"Macroregiunea patru"
"Y_GE15","RO41",2000,5,"Sud-Vest Oltenia"
"Y_GE15","RO42",2000,7.6,"Vest"
"Y_GE15","SE",2000,5.5,"Sweden"
"Y_GE15","SE1",2000,4.2,"Östra Sverige"
"Y_GE15","SE11",2000,3.2,"Stockholm"
"Y_GE15","SE12",2000,5.5,"Östra Mellansverige"
"Y_GE15","SE2",2000,5.7,"Södra Sverige"
"Y_GE15","SE21",2000,4.4,"Småland med öarna"
"Y_GE15","SE22",2000,7.3,"Sydsverige"
"Y_GE15","SE23",2000,5.2,"Västsverige"
"Y_GE15","SE3",2000,7.6,"Norra Sverige"
"Y_GE15","SE31",2000,6.7,"Norra Mellansverige"
"Y_GE15","SE32",2000,7.6,"Mellersta Norrland"
"Y_GE15","SE33",2000,9,"Övre Norrland"
"Y_GE15","SI",2000,6.9,"Slovenia"
"Y_GE15","SI0",2000,6.9,"Slovenija"
"Y_GE15","SK",2000,19.1,"Slovakia"
"Y_GE15","SK0",2000,19.1,"Slovensko"
"Y_GE15","SK01",2000,7.5,"Bratislavský kraj"
"Y_GE15","SK02",2000,17.6,"Západné Slovensko"
"Y_GE15","SK03",2000,21,"Stredné Slovensko"
"Y_GE15","SK04",2000,24.6,"Východné Slovensko"
"Y_GE15","UK",2000,5.6,"United Kingdom"
"Y_GE15","UKC",2000,9.1,"North East (UK)"
"Y_GE15","UKC1",2000,9,"Tees Valley and Durham"
"Y_GE15","UKC2",2000,9.2,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",2000,5.3,"North West (UK)"
"Y_GE15","UKD1",2000,5.1,"Cumbria"
"Y_GE15","UKD3",2000,5.1,"Greater Manchester"
"Y_GE15","UKD4",2000,4.5,"Lancashire"
"Y_GE15","UKE",2000,6,"Yorkshire and The Humber"
"Y_GE15","UKE1",2000,6.7,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",2000,4.9,"North Yorkshire"
"Y_GE15","UKE3",2000,6.9,"South Yorkshire"
"Y_GE15","UKE4",2000,5.6,"West Yorkshire"
"Y_GE15","UKF",2000,5.1,"East Midlands (UK)"
"Y_GE15","UKF1",2000,5.7,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",2000,4.7,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",2000,4.5,"Lincolnshire"
"Y_GE15","UKG",2000,6.3,"West Midlands (UK)"
"Y_GE15","UKG1",2000,4.2,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",2000,4.9,"Shropshire and Staffordshire"
"Y_GE15","UKG3",2000,8.2,"West Midlands"
"Y_GE15","UKH",2000,3.6,"East of England"
"Y_GE15","UKH1",2000,4.2,"East Anglia"
"Y_GE15","UKH2",2000,3.1,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",2000,3.4,"Essex"
"Y_GE15","UKI",2000,7.2,"London"
"Y_GE15","UKI1",2000,9.4,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",2000,5.7,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",2000,3.4,"South East (UK)"
"Y_GE15","UKJ1",2000,2.2,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",2000,3.1,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",2000,3.8,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",2000,5.1,"Kent"
"Y_GE15","UKK",2000,4.1,"South West (UK)"
"Y_GE15","UKK1",2000,3.2,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",2000,4.4,"Dorset and Somerset"
"Y_GE15","UKK3",2000,6.6,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",2000,4.9,"Devon"
"Y_GE15","UKL",2000,6.1,"Wales"
"Y_GE15","UKL1",2000,7,"West Wales and The Valleys"
"Y_GE15","UKL2",2000,4.9,"East Wales"
"Y_GE15","UKM",2000,7.6,"Scotland"
"Y_GE15","UKM2",2000,6.9,"Eastern Scotland"
"Y_GE15","UKM3",2000,9.1,"South Western Scotland"
"Y_GE15","UKM5",2000,NA,"North Eastern Scotland"
"Y_GE15","UKM6",2000,7.9,"Highlands and Islands"
"Y_GE15","UKN",2000,6.9,"Northern Ireland (UK)"
"Y_GE15","UKN0",2000,6.9,"Northern Ireland (UK)"
"Y_GE25","AT",2000,4.4,"Austria"
"Y_GE25","AT1",2000,5.7,"Ostösterreich"
"Y_GE25","AT11",2000,4.8,"Burgenland (AT)"
"Y_GE25","AT12",2000,4,"Niederösterreich"
"Y_GE25","AT13",2000,7.3,"Wien"
"Y_GE25","AT2",2000,4,"Südösterreich"
"Y_GE25","AT21",2000,4.2,"Kärnten"
"Y_GE25","AT22",2000,4,"Steiermark"
"Y_GE25","AT3",2000,3.2,"Westösterreich"
"Y_GE25","AT31",2000,3.6,"Oberösterreich"
"Y_GE25","AT32",2000,2.9,"Salzburg"
"Y_GE25","AT33",2000,2.8,"Tirol"
"Y_GE25","AT34",2000,NA,"Vorarlberg"
"Y_GE25","BE",2000,5.6,"Belgium"
"Y_GE25","BE1",2000,13.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",2000,13.1,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",2000,3,"Vlaams Gewest"
"Y_GE25","BE21",2000,3.6,"Prov. Antwerpen"
"Y_GE25","BE22",2000,4.3,"Prov. Limburg (BE)"
"Y_GE25","BE23",2000,2.6,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",2000,2.3,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",2000,2.6,"Prov. West-Vlaanderen"
"Y_GE25","BE3",2000,8.3,"Région wallonne"
"Y_GE25","BE31",2000,5.7,"Prov. Brabant Wallon"
"Y_GE25","BE32",2000,10.1,"Prov. Hainaut"
"Y_GE25","BE33",2000,7.7,"Prov. Liège"
"Y_GE25","BE34",2000,NA,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",2000,9,"Prov. Namur"
"Y_GE25","BG",2000,14.3,"Bulgaria"
"Y_GE25","BG41",2000,9.9,"Yugozapaden"
"Y_GE25","CH",2000,2.3,"Switzerland"
"Y_GE25","CH0",2000,2.3,"Schweiz/Suisse/Svizzera"
"Y_GE25","CY",2000,4.3,"Cyprus"
"Y_GE25","CY0",2000,4.3,"Kypros"
"Y_GE25","CY00",2000,4.3,"Kypros"
"Y_GE25","CZ",2000,7.5,"Czech Republic"
"Y_GE25","CZ0",2000,7.5,"Ceská republika"
"Y_GE25","CZ01",2000,3.2,"Praha"
"Y_GE25","CZ02",2000,6.9,"Strední Cechy"
"Y_GE25","CZ03",2000,5.2,"Jihozápad"
"Y_GE25","CZ04",2000,13.2,"Severozápad"
"Y_GE25","CZ05",2000,5.7,"Severovýchod"
"Y_GE25","CZ06",2000,6.3,"Jihovýchod"
"Y_GE25","CZ07",2000,9.5,"Strední Morava"
"Y_GE25","CZ08",2000,11.7,"Moravskoslezsko"
"Y_GE25","DE",2000,7.8,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",2000,3.9,"Baden-Württemberg"
"Y_GE25","DE11",2000,3.8,"Stuttgart"
"Y_GE25","DE12",2000,4.4,"Karlsruhe"
"Y_GE25","DE13",2000,4.1,"Freiburg"
"Y_GE25","DE14",2000,3.4,"Tübingen"
"Y_GE25","DE2",2000,3.9,"Bayern"
"Y_GE25","DE21",2000,2.9,"Oberbayern"
"Y_GE25","DE22",2000,3.3,"Niederbayern"
"Y_GE25","DE23",2000,4.7,"Oberpfalz"
"Y_GE25","DE24",2000,4.6,"Oberfranken"
"Y_GE25","DE25",2000,5.7,"Mittelfranken"
"Y_GE25","DE26",2000,4.2,"Unterfranken"
"Y_GE25","DE27",2000,3.8,"Schwaben"
"Y_GE25","DE3",2000,14.3,"Berlin"
"Y_GE25","DE30",2000,14.3,"Berlin"
"Y_GE25","DE4",2000,16.1,"Brandenburg"
"Y_GE25","DE40",2000,16.1,"Brandenburg"
"Y_GE25","DE5",2000,9.9,"Bremen"
"Y_GE25","DE50",2000,9.9,"Bremen"
"Y_GE25","DE6",2000,7.7,"Hamburg"
"Y_GE25","DE60",2000,7.7,"Hamburg"
"Y_GE25","DE7",2000,5.6,"Hessen"
"Y_GE25","DE71",2000,5.1,"Darmstadt"
"Y_GE25","DE72",2000,6.2,"Gießen"
"Y_GE25","DE73",2000,7,"Kassel"
"Y_GE25","DE8",2000,17.1,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",2000,17.1,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",2000,6.2,"Niedersachsen"
"Y_GE25","DE91",2000,6.9,"Braunschweig"
"Y_GE25","DE92",2000,7.2,"Hannover"
"Y_GE25","DE93",2000,5.9,"Lüneburg"
"Y_GE25","DE94",2000,5.2,"Weser-Ems"
"Y_GE25","DEA",2000,6.3,"Nordrhein-Westfalen"
"Y_GE25","DEA1",2000,6.5,"Düsseldorf"
"Y_GE25","DEA2",2000,5.8,"Köln"
"Y_GE25","DEA3",2000,5.3,"Münster"
"Y_GE25","DEA4",2000,5.6,"Detmold"
"Y_GE25","DEA5",2000,7.5,"Arnsberg"
"Y_GE25","DEB",2000,5.5,"Rheinland-Pfalz"
"Y_GE25","DEC",2000,6.9,"Saarland"
"Y_GE25","DEC0",2000,6.9,"Saarland"
"Y_GE25","DED",2000,16.5,"Sachsen"
"Y_GE25","DED2",2000,16.5,"Dresden"
"Y_GE25","DEE",2000,21.2,"Sachsen-Anhalt"
"Y_GE25","DEE0",2000,21.2,"Sachsen-Anhalt"
"Y_GE25","DEF",2000,6.3,"Schleswig-Holstein"
"Y_GE25","DEF0",2000,6.3,"Schleswig-Holstein"
"Y_GE25","DEG",2000,14,"Thüringen"
"Y_GE25","DEG0",2000,14,"Thüringen"
"Y_GE25","DK",2000,4.1,"Denmark"
"Y_GE25","DK0",2000,4.1,"Danmark"
"Y_GE25","EA17",2000,8.1,"Euro area (17 countries)"
"Y_GE25","EA18",2000,8.2,"Euro area (18 countries)"
"Y_GE25","EA19",2000,8.2,"Euro area (19 countries)"
"Y_GE25","EE",2000,12.4,"Estonia"
"Y_GE25","EE0",2000,12.4,"Eesti"
"Y_GE25","EE00",2000,12.4,"Eesti"
"Y_GE25","EL",2000,8.8,"Greece"
"Y_GE25","EL1",2000,8.9,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",2000,7.2,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",2000,8.5,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",2000,11.5,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",2000,10.3,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",2000,7.8,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",2000,8.9,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",2000,4.9,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",2000,7,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",2000,10,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",2000,7.1,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",2000,10,"Attiki"
"Y_GE25","EL30",2000,10,"Attiki"
"Y_GE25","EL4",2000,6,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",2000,6.1,"Voreio Aigaio"
"Y_GE25","EL42",2000,8.5,"Notio Aigaio"
"Y_GE25","EL43",2000,4.8,"Kriti"
"Y_GE25","ES",2000,11.9,"Spain"
"Y_GE25","ES1",2000,13.1,"Noroeste (ES)"
"Y_GE25","ES11",2000,12.8,"Galicia"
"Y_GE25","ES12",2000,15,"Principado de Asturias"
"Y_GE25","ES13",2000,11,"Cantabria"
"Y_GE25","ES2",2000,7.9,"Noreste (ES)"
"Y_GE25","ES21",2000,10.4,"País Vasco"
"Y_GE25","ES22",2000,3.4,"Comunidad Foral de Navarra"
"Y_GE25","ES23",2000,6.2,"La Rioja"
"Y_GE25","ES24",2000,5.7,"Aragón"
"Y_GE25","ES3",2000,10,"Comunidad de Madrid"
"Y_GE25","ES30",2000,10,"Comunidad de Madrid"
"Y_GE25","ES4",2000,13.5,"Centro (ES)"
"Y_GE25","ES41",2000,11.7,"Castilla y León"
"Y_GE25","ES42",2000,10.8,"Castilla-la Mancha"
"Y_GE25","ES43",2000,22.4,"Extremadura"
"Y_GE25","ES5",2000,7.8,"Este (ES)"
"Y_GE25","ES51",2000,7.1,"Cataluña"
"Y_GE25","ES52",2000,9.8,"Comunidad Valenciana"
"Y_GE25","ES53",2000,4.4,"Illes Balears"
"Y_GE25","ES6",2000,20,"Sur (ES)"
"Y_GE25","ES61",2000,21.8,"Andalucía"
"Y_GE25","ES62",2000,9,"Región de Murcia"
"Y_GE25","ES63",2000,21.8,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",2000,18.3,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",2000,12.2,"Canarias (ES)"
"Y_GE25","ES70",2000,12.2,"Canarias (ES)"
"Y_GE25","EU15",2000,7.3,"European Union (15 countries)"
"Y_GE25","EU27",2000,7.9,"European Union (27 countries)"
"Y_GE25","FI",2000,8,"Finland"
"Y_GE25","FI1",2000,8.1,"Manner-Suomi"
"Y_GE25","FI19",2000,8.2,"Länsi-Suomi"
"Y_GE25","FI2",2000,NA,"Åland"
"Y_GE25","FI20",2000,NA,"Åland"
"Y_GE25","FR",2000,9.1,"France"
"Y_GE25","FR1",2000,8.1,"Île de France"
"Y_GE25","FR10",2000,8.1,"Île de France"
"Y_GE25","FR2",2000,8.8,"Bassin Parisien"
"Y_GE25","FR21",2000,9.8,"Champagne-Ardenne"
"Y_GE25","FR22",2000,9.9,"Picardie"
"Y_GE25","FR23",2000,10,"Haute-Normandie"
"Y_GE25","FR24",2000,7.3,"Centre (FR)"
"Y_GE25","FR25",2000,7.4,"Basse-Normandie"
"Y_GE25","FR26",2000,8.5,"Bourgogne"
"Y_GE25","FR3",2000,13.8,"Nord - Pas-de-Calais"
"Y_GE25","FR30",2000,13.8,"Nord - Pas-de-Calais"
"Y_GE25","FR4",2000,7.3,"Est (FR)"
"Y_GE25","FR41",2000,8.7,"Lorraine"
"Y_GE25","FR42",2000,5.7,"Alsace"
"Y_GE25","FR43",2000,6.9,"Franche-Comté"
"Y_GE25","FR5",2000,7.6,"Ouest (FR)"
"Y_GE25","FR51",2000,8.6,"Pays de la Loire"
"Y_GE25","FR52",2000,6.4,"Bretagne"
"Y_GE25","FR53",2000,7.4,"Poitou-Charentes"
"Y_GE25","FR6",2000,9.1,"Sud-Ouest (FR)"
"Y_GE25","FR61",2000,9.7,"Aquitaine"
"Y_GE25","FR62",2000,9,"Midi-Pyrénées"
"Y_GE25","FR63",2000,6.9,"Limousin"
"Y_GE25","FR7",2000,7.5,"Centre-Est (FR)"
"Y_GE25","FR71",2000,7.1,"Rhône-Alpes"
"Y_GE25","FR72",2000,8.9,"Auvergne"
"Y_GE25","FR8",2000,14.1,"Méditerranée"
"Y_GE25","FR81",2000,14.6,"Languedoc-Roussillon"
"Y_GE25","FR82",2000,13.6,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",2000,NA,"Corse"
"Y_GE25","HU",2000,5.6,"Hungary"
"Y_GE25","HU1",2000,4.5,"Közép-Magyarország"
"Y_GE25","HU10",2000,4.5,"Közép-Magyarország"
"Y_GE25","HU2",2000,5.1,"Dunántúl"
"Y_GE25","HU21",2000,4.7,"Közép-Dunántúl"
"Y_GE25","HU22",2000,3.7,"Nyugat-Dunántúl"
"Y_GE25","HU23",2000,7.2,"Dél-Dunántúl"
"Y_GE25","HU3",2000,7,"Alföld és Észak"
"Y_GE25","HU31",2000,8.2,"Észak-Magyarország"
"Y_GE25","HU32",2000,8.5,"Észak-Alföld"
"Y_GE25","HU33",2000,4.6,"Dél-Alföld"
"Y_GE25","IE",2000,3.8,"Ireland"
"Y_GE25","IE0",2000,3.8,"Éire/Ireland"
"Y_GE25","IE01",2000,4.8,"Border, Midland and Western"
"Y_GE25","IE02",2000,3.5,"Southern and Eastern"
"Y_GE25","IS",2000,1.4,"Iceland"
"Y_GE25","IS0",2000,1.4,"Ísland"
"Y_GE25","IS00",2000,1.4,"Ísland"
"Y_GE25","IT",2000,8.3,"Italy"
"Y_GE25","ITC",2000,4.2,"Nord-Ovest"
"Y_GE25","ITC1",2000,5,"Piemonte"
"Y_GE25","ITC2",2000,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",2000,7.1,"Liguria"
"Y_GE25","ITC4",2000,3.4,"Lombardia"
"Y_GE25","ITF",2000,15.1,"Sud"
"Y_GE25","ITF1",2000,5.8,"Abruzzo"
"Y_GE25","ITF2",2000,9.5,"Molise"
"Y_GE25","ITF3",2000,17.2,"Campania"
"Y_GE25","ITF4",2000,12.6,"Puglia"
"Y_GE25","ITF5",2000,14.3,"Basilicata"
"Y_GE25","ITF6",2000,22.1,"Calabria"
"Y_GE25","ITG",2000,17.8,"Isole"
"Y_GE25","ITG1",2000,18.5,"Sicilia"
"Y_GE25","ITG2",2000,16,"Sardegna"
"Y_GE25","ITH",2000,3.6,"Nord-Est"
"Y_GE25","ITH1",2000,2,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",2000,3,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",2000,3.5,"Veneto"
"Y_GE25","ITH4",2000,3.8,"Friuli-Venezia Giulia"
"Y_GE25","ITI",2000,7,"Centro (IT)"
"Y_GE25","ITI1",2000,5.5,"Toscana"
"Y_GE25","ITI2",2000,4.8,"Umbria"
"Y_GE25","ITI4",2000,9.2,"Lazio"
"Y_GE25","LT",2000,14.4,"Lithuania"
"Y_GE25","LT0",2000,14.4,"Lietuva"
"Y_GE25","LT00",2000,14.4,"Lietuva"
"Y_GE25","LU",2000,2,"Luxembourg"
"Y_GE25","LU0",2000,2,"Luxembourg"
"Y_GE25","LU00",2000,2,"Luxembourg"
"Y_GE25","LV",2000,13.3,"Latvia"
"Y_GE25","LV0",2000,13.3,"Latvija"
"Y_GE25","LV00",2000,13.3,"Latvija"
"Y_GE25","MT",2000,4.7,"Malta"
"Y_GE25","MT0",2000,4.7,"Malta"
"Y_GE25","MT00",2000,4.7,"Malta"
"Y_GE25","NL",2000,2.2,"Netherlands"
"Y_GE25","NL1",2000,3.6,"Noord-Nederland"
"Y_GE25","NL11",2000,3.8,"Groningen"
"Y_GE25","NL12",2000,3.8,"Friesland (NL)"
"Y_GE25","NL13",2000,3.1,"Drenthe"
"Y_GE25","NL2",2000,2.2,"Oost-Nederland"
"Y_GE25","NL21",2000,1.9,"Overijssel"
"Y_GE25","NL22",2000,2,"Gelderland"
"Y_GE25","NL23",2000,4,"Flevoland"
"Y_GE25","NL3",2000,2.1,"West-Nederland"
"Y_GE25","NL31",2000,1.3,"Utrecht"
"Y_GE25","NL32",2000,2.5,"Noord-Holland"
"Y_GE25","NL33",2000,2,"Zuid-Holland"
"Y_GE25","NL34",2000,2.9,"Zeeland"
"Y_GE25","NL4",2000,1.9,"Zuid-Nederland"
"Y_GE25","NL41",2000,1.8,"Noord-Brabant"
"Y_GE25","NL42",2000,2.3,"Limburg (NL)"
"Y_GE25","NO",2000,2.2,"Norway"
"Y_GE25","NO0",2000,2.2,"Norge"
"Y_GE25","NO01",2000,1.8,"Oslo og Akershus"
"Y_GE25","NO02",2000,2.1,"Hedmark og Oppland"
"Y_GE25","NO03",2000,1.9,"Sør-Østlandet"
"Y_GE25","NO04",2000,2.9,"Agder og Rogaland"
"Y_GE25","NO05",2000,2.4,"Vestlandet"
"Y_GE25","NO06",2000,2.1,"Trøndelag"
"Y_GE25","NO07",2000,2.4,"Nord-Norge"
"Y_GE25","PL",2000,13.6,"Poland"
"Y_GE25","PL1",2000,11.5,"Region Centralny"
"Y_GE25","PL11",2000,12.9,"Lódzkie"
"Y_GE25","PL12",2000,10.7,"Mazowieckie"
"Y_GE25","PL2",2000,13,"Region Poludniowy"
"Y_GE25","PL21",2000,9.3,"Malopolskie"
"Y_GE25","PL22",2000,16.5,"Slaskie"
"Y_GE25","PL3",2000,12.1,"Region Wschodni"
"Y_GE25","PL31",2000,11,"Lubelskie"
"Y_GE25","PL32",2000,11.5,"Podkarpackie"
"Y_GE25","PL33",2000,13.7,"Swietokrzyskie"
"Y_GE25","PL34",2000,13.9,"Podlaskie"
"Y_GE25","PL4",2000,13.9,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",2000,10.9,"Wielkopolskie"
"Y_GE25","PL42",2000,17.2,"Zachodniopomorskie"
"Y_GE25","PL43",2000,19.3,"Lubuskie"
"Y_GE25","PL5",2000,17.8,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",2000,19.9,"Dolnoslaskie"
"Y_GE25","PL52",2000,12.5,"Opolskie"
"Y_GE25","PL6",2000,16.3,"Region Pólnocny"
"Y_GE25","PL61",2000,15.5,"Kujawsko-Pomorskie"
"Y_GE25","PL62",2000,19.1,"Warminsko-Mazurskie"
"Y_GE25","PL63",2000,14.8,"Pomorskie"
"Y_GE25","PT",2000,3.2,"Portugal"
"Y_GE25","PT1",2000,3.2,"Continente"
"Y_GE25","PT11",2000,3.3,"Norte"
"Y_GE25","PT15",2000,NA,"Algarve"
"Y_GE25","PT16",2000,1.2,"Centro (PT)"
"Y_GE25","PT17",2000,4.7,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",2000,4.9,"Alentejo"
"Y_GE25","PT2",2000,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",2000,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",2000,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",2000,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",2000,5.4,"Romania"
"Y_GE25","RO1",2000,5.8,"Macroregiunea unu"
"Y_GE25","RO11",2000,5.6,"Nord-Vest"
"Y_GE25","RO12",2000,6,"Centru"
"Y_GE25","RO2",2000,6.2,"Macroregiunea doi"
"Y_GE25","RO21",2000,5.4,"Nord-Est"
"Y_GE25","RO22",2000,7.3,"Sud-Est"
"Y_GE25","RO3",2000,4.8,"Macroregiunea trei"
"Y_GE25","RO31",2000,4.6,"Sud - Muntenia"
"Y_GE25","RO32",2000,5.1,"Bucuresti - Ilfov"
"Y_GE25","RO4",2000,4.6,"Macroregiunea patru"
"Y_GE25","RO41",2000,3.9,"Sud-Vest Oltenia"
"Y_GE25","RO42",2000,5.7,"Vest"
"Y_GE25","SE",2000,5,"Sweden"
"Y_GE25","SE1",2000,3.7,"Östra Sverige"
"Y_GE25","SE11",2000,2.9,"Stockholm"
"Y_GE25","SE12",2000,4.9,"Östra Mellansverige"
"Y_GE25","SE2",2000,5.3,"Södra Sverige"
"Y_GE25","SE21",2000,4.3,"Småland med öarna"
"Y_GE25","SE22",2000,6.4,"Sydsverige"
"Y_GE25","SE23",2000,5.1,"Västsverige"
"Y_GE25","SE3",2000,7.1,"Norra Sverige"
"Y_GE25","SE31",2000,5.9,"Norra Mellansverige"
"Y_GE25","SE32",2000,7.4,"Mellersta Norrland"
"Y_GE25","SE33",2000,8.8,"Övre Norrland"
"Y_GE25","SI",2000,5.7,"Slovenia"
"Y_GE25","SI0",2000,5.7,"Slovenija"
"Y_GE25","SK",2000,15.7,"Slovakia"
"Y_GE25","SK0",2000,15.7,"Slovensko"
"Y_GE25","SK01",2000,5.9,"Bratislavský kraj"
"Y_GE25","SK02",2000,14.8,"Západné Slovensko"
"Y_GE25","SK03",2000,17.7,"Stredné Slovensko"
"Y_GE25","SK04",2000,20.1,"Východné Slovensko"
"Y_GE25","UK",2000,4.4,"United Kingdom"
"Y_GE25","UKC",2000,7,"North East (UK)"
"Y_GE25","UKC1",2000,6.4,"Tees Valley and Durham"
"Y_GE25","UKC2",2000,7.5,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",2000,4.5,"North West (UK)"
"Y_GE25","UKD1",2000,NA,"Cumbria"
"Y_GE25","UKD3",2000,4.1,"Greater Manchester"
"Y_GE25","UKD4",2000,3.7,"Lancashire"
"Y_GE25","UKE",2000,4.7,"Yorkshire and The Humber"
"Y_GE25","UKE1",2000,5.5,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",2000,3.3,"North Yorkshire"
"Y_GE25","UKE3",2000,5.4,"South Yorkshire"
"Y_GE25","UKE4",2000,4.5,"West Yorkshire"
"Y_GE25","UKF",2000,3.8,"East Midlands (UK)"
"Y_GE25","UKF1",2000,4.3,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",2000,3.6,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",2000,NA,"Lincolnshire"
"Y_GE25","UKG",2000,4.9,"West Midlands (UK)"
"Y_GE25","UKG1",2000,3.7,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",2000,4.1,"Shropshire and Staffordshire"
"Y_GE25","UKG3",2000,6.1,"West Midlands"
"Y_GE25","UKH",2000,2.8,"East of England"
"Y_GE25","UKH1",2000,3.5,"East Anglia"
"Y_GE25","UKH2",2000,2.2,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",2000,2.6,"Essex"
"Y_GE25","UKI",2000,5.8,"London"
"Y_GE25","UKI1",2000,7.8,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",2000,4.5,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",2000,2.8,"South East (UK)"
"Y_GE25","UKJ1",2000,1.7,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",2000,2.7,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",2000,3,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",2000,4.2,"Kent"
"Y_GE25","UKK",2000,3.3,"South West (UK)"
"Y_GE25","UKK1",2000,2.4,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",2000,3.9,"Dorset and Somerset"
"Y_GE25","UKK3",2000,5.7,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",2000,3.8,"Devon"
"Y_GE25","UKL",2000,4.7,"Wales"
"Y_GE25","UKL1",2000,5.4,"West Wales and The Valleys"
"Y_GE25","UKL2",2000,3.6,"East Wales"
"Y_GE25","UKM",2000,6.1,"Scotland"
"Y_GE25","UKM2",2000,5.3,"Eastern Scotland"
"Y_GE25","UKM3",2000,7.4,"South Western Scotland"
"Y_GE25","UKM5",2000,NA,"North Eastern Scotland"
"Y_GE25","UKM6",2000,6.7,"Highlands and Islands"
"Y_GE25","UKN",2000,6,"Northern Ireland (UK)"
"Y_GE25","UKN0",2000,6,"Northern Ireland (UK)"
"Y15-24","AT",1999,5.9,"Austria"
"Y15-24","AT1",1999,6.1,"Ostösterreich"
"Y15-24","AT11",1999,NA,"Burgenland (AT)"
"Y15-24","AT12",1999,4.4,"Niederösterreich"
"Y15-24","AT13",1999,7.9,"Wien"
"Y15-24","AT2",1999,5.2,"Südösterreich"
"Y15-24","AT21",1999,NA,"Kärnten"
"Y15-24","AT22",1999,5.4,"Steiermark"
"Y15-24","AT3",1999,6.2,"Westösterreich"
"Y15-24","AT31",1999,7.2,"Oberösterreich"
"Y15-24","AT32",1999,NA,"Salzburg"
"Y15-24","AT33",1999,NA,"Tirol"
"Y15-24","AT34",1999,NA,"Vorarlberg"
"Y15-24","BE",1999,22.6,"Belgium"
"Y15-24","BE1",1999,37,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE10",1999,37,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y15-24","BE2",1999,15.6,"Vlaams Gewest"
"Y15-24","BE21",1999,18.2,"Prov. Antwerpen"
"Y15-24","BE22",1999,15.9,"Prov. Limburg (BE)"
"Y15-24","BE23",1999,16.7,"Prov. Oost-Vlaanderen"
"Y15-24","BE24",1999,14.7,"Prov. Vlaams-Brabant"
"Y15-24","BE25",1999,11.4,"Prov. West-Vlaanderen"
"Y15-24","BE3",1999,32.3,"Région wallonne"
"Y15-24","BE31",1999,NA,"Prov. Brabant Wallon"
"Y15-24","BE32",1999,37,"Prov. Hainaut"
"Y15-24","BE33",1999,31.7,"Prov. Liège"
"Y15-24","BE34",1999,NA,"Prov. Luxembourg (BE)"
"Y15-24","BE35",1999,34.5,"Prov. Namur"
"Y15-24","CH",1999,6.2,"Switzerland"
"Y15-24","CH0",1999,6.2,"Schweiz/Suisse/Svizzera"
"Y15-24","CZ",1999,16.6,"Czech Republic"
"Y15-24","CZ0",1999,16.6,"Ceská republika"
"Y15-24","CZ01",1999,9.1,"Praha"
"Y15-24","CZ02",1999,13.4,"Strední Cechy"
"Y15-24","CZ03",1999,10.9,"Jihozápad"
"Y15-24","CZ04",1999,23.1,"Severozápad"
"Y15-24","CZ05",1999,15.2,"Severovýchod"
"Y15-24","CZ06",1999,15.1,"Jihovýchod"
"Y15-24","CZ07",1999,18.7,"Strední Morava"
"Y15-24","CZ08",1999,26,"Moravskoslezsko"
"Y15-24","DE",1999,8.9,"Germany (until 1990 former territory of the FRG)"
"Y15-24","DE1",1999,5.1,"Baden-Württemberg"
"Y15-24","DE11",1999,4.2,"Stuttgart"
"Y15-24","DE12",1999,5.2,"Karlsruhe"
"Y15-24","DE13",1999,6.7,"Freiburg"
"Y15-24","DE14",1999,5.3,"Tübingen"
"Y15-24","DE2",1999,6.1,"Bayern"
"Y15-24","DE21",1999,4.9,"Oberbayern"
"Y15-24","DE22",1999,NA,"Niederbayern"
"Y15-24","DE23",1999,NA,"Oberpfalz"
"Y15-24","DE24",1999,7.9,"Oberfranken"
"Y15-24","DE25",1999,8.3,"Mittelfranken"
"Y15-24","DE26",1999,9.4,"Unterfranken"
"Y15-24","DE27",1999,5.4,"Schwaben"
"Y15-24","DE3",1999,16.6,"Berlin"
"Y15-24","DE30",1999,16.6,"Berlin"
"Y15-24","DE4",1999,13.9,"Brandenburg"
"Y15-24","DE40",1999,13.9,"Brandenburg"
"Y15-24","DE5",1999,NA,"Bremen"
"Y15-24","DE50",1999,NA,"Bremen"
"Y15-24","DE6",1999,10,"Hamburg"
"Y15-24","DE60",1999,10,"Hamburg"
"Y15-24","DE7",1999,9,"Hessen"
"Y15-24","DE71",1999,8.6,"Darmstadt"
"Y15-24","DE72",1999,10.7,"Gießen"
"Y15-24","DE73",1999,8.6,"Kassel"
"Y15-24","DE8",1999,11,"Mecklenburg-Vorpommern"
"Y15-24","DE80",1999,11,"Mecklenburg-Vorpommern"
"Y15-24","DE9",1999,8.7,"Niedersachsen"
"Y15-24","DE91",1999,12,"Braunschweig"
"Y15-24","DE92",1999,6.8,"Hannover"
"Y15-24","DE93",1999,8.7,"Lüneburg"
"Y15-24","DE94",1999,7.8,"Weser-Ems"
"Y15-24","DEA",1999,9.6,"Nordrhein-Westfalen"
"Y15-24","DEA1",1999,11,"Düsseldorf"
"Y15-24","DEA2",1999,7.7,"Köln"
"Y15-24","DEA3",1999,11.3,"Münster"
"Y15-24","DEA4",1999,6.7,"Detmold"
"Y15-24","DEA5",1999,10.5,"Arnsberg"
"Y15-24","DEB",1999,7.2,"Rheinland-Pfalz"
"Y15-24","DEB1",1999,10.4,"Koblenz"
"Y15-24","DEB2",1999,NA,"Trier"
"Y15-24","DEB3",1999,5.3,"Rheinhessen-Pfalz"
"Y15-24","DEC",1999,NA,"Saarland"
"Y15-24","DEC0",1999,NA,"Saarland"
"Y15-24","DED",1999,10.9,"Sachsen"
"Y15-24","DEE",1999,12.5,"Sachsen-Anhalt"
"Y15-24","DEE0",1999,12.5,"Sachsen-Anhalt"
"Y15-24","DEF",1999,10.1,"Schleswig-Holstein"
"Y15-24","DEF0",1999,10.1,"Schleswig-Holstein"
"Y15-24","DEG",1999,8.3,"Thüringen"
"Y15-24","DEG0",1999,8.3,"Thüringen"
"Y15-24","DK",1999,10,"Denmark"
"Y15-24","DK0",1999,10,"Danmark"
"Y15-24","EE",1999,22.1,"Estonia"
"Y15-24","EE0",1999,22.1,"Eesti"
"Y15-24","EE00",1999,22.1,"Eesti"
"Y15-24","EL",1999,31.4,"Greece"
"Y15-24","EL1",1999,31.9,"Voreia Ellada (NUTS 2010)"
"Y15-24","EL11",1999,30.8,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y15-24","EL12",1999,29.8,"Kentriki Makedonia (NUTS 2010)"
"Y15-24","EL13",1999,46.4,"Dytiki Makedonia (NUTS 2010)"
"Y15-24","EL14",1999,33.2,"Thessalia (NUTS 2010)"
"Y15-24","EL2",1999,34.1,"Kentriki Ellada (NUTS 2010)"
"Y15-24","EL21",1999,42,"Ipeiros (NUTS 2010)"
"Y15-24","EL22",1999,21.1,"Ionia Nisia (NUTS 2010)"
"Y15-24","EL23",1999,36.7,"Dytiki Ellada (NUTS 2010)"
"Y15-24","EL24",1999,37.9,"Sterea Ellada (NUTS 2010)"
"Y15-24","EL25",1999,27,"Peloponnisos (NUTS 2010)"
"Y15-24","EL3",1999,33,"Attiki"
"Y15-24","EL30",1999,33,"Attiki"
"Y15-24","EL4",1999,19.9,"Nisia Aigaiou, Kriti"
"Y15-24","EL41",1999,28.3,"Voreio Aigaio"
"Y15-24","EL42",1999,16,"Notio Aigaio"
"Y15-24","EL43",1999,20,"Kriti"
"Y15-24","ES",1999,29.1,"Spain"
"Y15-24","ES1",1999,34.6,"Noroeste (ES)"
"Y15-24","ES11",1999,31.8,"Galicia"
"Y15-24","ES12",1999,44.2,"Principado de Asturias"
"Y15-24","ES13",1999,31.7,"Cantabria"
"Y15-24","ES2",1999,22.8,"Noreste (ES)"
"Y15-24","ES21",1999,30,"País Vasco"
"Y15-24","ES22",1999,14.8,"Comunidad Foral de Navarra"
"Y15-24","ES23",1999,NA,"La Rioja"
"Y15-24","ES24",1999,16.4,"Aragón"
"Y15-24","ES3",1999,25,"Comunidad de Madrid"
"Y15-24","ES30",1999,25,"Comunidad de Madrid"
"Y15-24","ES4",1999,32.8,"Centro (ES)"
"Y15-24","ES41",1999,34.4,"Castilla y León"
"Y15-24","ES42",1999,26.3,"Castilla-la Mancha"
"Y15-24","ES43",1999,41.1,"Extremadura"
"Y15-24","ES5",1999,22,"Este (ES)"
"Y15-24","ES51",1999,20.6,"Cataluña"
"Y15-24","ES52",1999,25.9,"Comunidad Valenciana"
"Y15-24","ES53",1999,13.8,"Illes Balears"
"Y15-24","ES6",1999,39.2,"Sur (ES)"
"Y15-24","ES61",1999,41.3,"Andalucía"
"Y15-24","ES62",1999,25.7,"Región de Murcia"
"Y15-24","ES63",1999,48.7,"Ciudad Autónoma de Ceuta (ES)"
"Y15-24","ES64",1999,NA,"Ciudad Autónoma de Melilla (ES)"
"Y15-24","ES7",1999,28.7,"Canarias (ES)"
"Y15-24","ES70",1999,28.7,"Canarias (ES)"
"Y15-24","EU15",1999,18.2,"European Union (15 countries)"
"Y15-24","FI",1999,28.6,"Finland"
"Y15-24","FI1",1999,28.6,"Manner-Suomi"
"Y15-24","FI19",1999,30.2,"Länsi-Suomi"
"Y15-24","FR",1999,26.3,"France"
"Y15-24","FR1",1999,21.4,"Île de France"
"Y15-24","FR10",1999,21.4,"Île de France"
"Y15-24","FR2",1999,27.6,"Bassin Parisien"
"Y15-24","FR21",1999,30.3,"Champagne-Ardenne"
"Y15-24","FR22",1999,31,"Picardie"
"Y15-24","FR23",1999,35.9,"Haute-Normandie"
"Y15-24","FR24",1999,21.1,"Centre (FR)"
"Y15-24","FR25",1999,24.2,"Basse-Normandie"
"Y15-24","FR26",1999,23.2,"Bourgogne"
"Y15-24","FR3",1999,42.4,"Nord - Pas-de-Calais"
"Y15-24","FR30",1999,42.4,"Nord - Pas-de-Calais"
"Y15-24","FR4",1999,20.2,"Est (FR)"
"Y15-24","FR41",1999,23.7,"Lorraine"
"Y15-24","FR42",1999,16.5,"Alsace"
"Y15-24","FR43",1999,NA,"Franche-Comté"
"Y15-24","FR5",1999,25.3,"Ouest (FR)"
"Y15-24","FR51",1999,23.7,"Pays de la Loire"
"Y15-24","FR52",1999,25.4,"Bretagne"
"Y15-24","FR53",1999,29,"Poitou-Charentes"
"Y15-24","FR6",1999,27.6,"Sud-Ouest (FR)"
"Y15-24","FR61",1999,28.5,"Aquitaine"
"Y15-24","FR62",1999,26.8,"Midi-Pyrénées"
"Y15-24","FR63",1999,NA,"Limousin"
"Y15-24","FR7",1999,22.5,"Centre-Est (FR)"
"Y15-24","FR71",1999,21.1,"Rhône-Alpes"
"Y15-24","FR72",1999,30.2,"Auvergne"
"Y15-24","FR8",1999,30.7,"Méditerranée"
"Y15-24","FR81",1999,31.5,"Languedoc-Roussillon"
"Y15-24","FR82",1999,29.3,"Provence-Alpes-Côte d'Azur"
"Y15-24","FR83",1999,NA,"Corse"
"Y15-24","HU",1999,12.3,"Hungary"
"Y15-24","HU1",1999,8.4,"Közép-Magyarország"
"Y15-24","HU10",1999,8.4,"Közép-Magyarország"
"Y15-24","HU2",1999,10.7,"Dunántúl"
"Y15-24","HU21",1999,9.4,"Közép-Dunántúl"
"Y15-24","HU22",1999,6.5,"Nyugat-Dunántúl"
"Y15-24","HU23",1999,17.4,"Dél-Dunántúl"
"Y15-24","HU3",1999,16.2,"Alföld és Észak"
"Y15-24","HU31",1999,20.8,"Észak-Magyarország"
"Y15-24","HU32",1999,16.7,"Észak-Alföld"
"Y15-24","HU33",1999,11.8,"Dél-Alföld"
"Y15-24","IE",1999,8.6,"Ireland"
"Y15-24","IE0",1999,8.6,"Éire/Ireland"
"Y15-24","IE01",1999,10.3,"Border, Midland and Western"
"Y15-24","IE02",1999,8.1,"Southern and Eastern"
"Y15-24","IS",1999,4.3,"Iceland"
"Y15-24","IS0",1999,4.3,"Ísland"
"Y15-24","IS00",1999,4.3,"Ísland"
"Y15-24","IT",1999,32.9,"Italy"
"Y15-24","ITC",1999,17.6,"Nord-Ovest"
"Y15-24","ITC1",1999,22.4,"Piemonte"
"Y15-24","ITC2",1999,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y15-24","ITC3",1999,31.2,"Liguria"
"Y15-24","ITC4",1999,13.7,"Lombardia"
"Y15-24","ITF",1999,55.1,"Sud"
"Y15-24","ITF1",1999,31.6,"Abruzzo"
"Y15-24","ITF2",1999,50.4,"Molise"
"Y15-24","ITF3",1999,60.9,"Campania"
"Y15-24","ITF4",1999,49,"Puglia"
"Y15-24","ITF5",1999,52.8,"Basilicata"
"Y15-24","ITF6",1999,65.2,"Calabria"
"Y15-24","ITG",1999,59.4,"Isole"
"Y15-24","ITG1",1999,60.2,"Sicilia"
"Y15-24","ITG2",1999,56.7,"Sardegna"
"Y15-24","ITH",1999,11.6,"Nord-Est"
"Y15-24","ITH1",1999,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y15-24","ITH2",1999,NA,"Provincia Autonoma di Trento"
"Y15-24","ITH3",1999,11.5,"Veneto"
"Y15-24","ITH4",1999,12.1,"Friuli-Venezia Giulia"
"Y15-24","ITI",1999,31.4,"Centro (IT)"
"Y15-24","ITI1",1999,20.8,"Toscana"
"Y15-24","ITI2",1999,19.9,"Umbria"
"Y15-24","ITI4",1999,46.9,"Lazio"
"Y15-24","LT",1999,25.5,"Lithuania"
"Y15-24","LT0",1999,25.5,"Lietuva"
"Y15-24","LT00",1999,25.5,"Lietuva"
"Y15-24","LU",1999,6.8,"Luxembourg"
"Y15-24","LU0",1999,6.8,"Luxembourg"
"Y15-24","LU00",1999,6.8,"Luxembourg"
"Y15-24","LV",1999,23.5,"Latvia"
"Y15-24","LV0",1999,23.5,"Latvija"
"Y15-24","LV00",1999,23.5,"Latvija"
"Y15-24","NL",1999,7.4,"Netherlands"
"Y15-24","NL1",1999,12.3,"Noord-Nederland"
"Y15-24","NL11",1999,13.2,"Groningen"
"Y15-24","NL12",1999,9.5,"Friesland (NL)"
"Y15-24","NL13",1999,15.8,"Drenthe"
"Y15-24","NL2",1999,7.2,"Oost-Nederland"
"Y15-24","NL21",1999,7.1,"Overijssel"
"Y15-24","NL22",1999,7.4,"Gelderland"
"Y15-24","NL23",1999,6.3,"Flevoland"
"Y15-24","NL3",1999,6.9,"West-Nederland"
"Y15-24","NL31",1999,2.6,"Utrecht"
"Y15-24","NL32",1999,7.2,"Noord-Holland"
"Y15-24","NL33",1999,7.9,"Zuid-Holland"
"Y15-24","NL34",1999,9.6,"Zeeland"
"Y15-24","NL4",1999,6.1,"Zuid-Nederland"
"Y15-24","NL41",1999,5.8,"Noord-Brabant"
"Y15-24","NL42",1999,6.8,"Limburg (NL)"
"Y15-24","NO",1999,12.3,"Norway"
"Y15-24","NO0",1999,12.3,"Norge"
"Y15-24","NO01",1999,10.1,"Oslo og Akershus"
"Y15-24","NO02",1999,18,"Hedmark og Oppland"
"Y15-24","NO03",1999,12.1,"Sør-Østlandet"
"Y15-24","NO04",1999,9.5,"Agder og Rogaland"
"Y15-24","NO05",1999,11.4,"Vestlandet"
"Y15-24","NO06",1999,15.1,"Trøndelag"
"Y15-24","NO07",1999,17.4,"Nord-Norge"
"Y15-24","PL",1999,29.6,"Poland"
"Y15-24","PL1",1999,23.8,"Region Centralny"
"Y15-24","PL11",1999,26,"Lódzkie"
"Y15-24","PL12",1999,22.6,"Mazowieckie"
"Y15-24","PL2",1999,26.3,"Region Poludniowy"
"Y15-24","PL21",1999,30.9,"Malopolskie"
"Y15-24","PL22",1999,23,"Slaskie"
"Y15-24","PL3",1999,34.2,"Region Wschodni"
"Y15-24","PL31",1999,31.9,"Lubelskie"
"Y15-24","PL32",1999,43.3,"Podkarpackie"
"Y15-24","PL33",1999,33.4,"Swietokrzyskie"
"Y15-24","PL34",1999,26.5,"Podlaskie"
"Y15-24","PL4",1999,32.9,"Region Pólnocno-Zachodni"
"Y15-24","PL41",1999,24.9,"Wielkopolskie"
"Y15-24","PL42",1999,53.1,"Zachodniopomorskie"
"Y15-24","PL43",1999,26.1,"Lubuskie"
"Y15-24","PL5",1999,34.6,"Region Poludniowo-Zachodni"
"Y15-24","PL51",1999,35.5,"Dolnoslaskie"
"Y15-24","PL52",1999,32.3,"Opolskie"
"Y15-24","PL6",1999,29.4,"Region Pólnocny"
"Y15-24","PL61",1999,31,"Kujawsko-Pomorskie"
"Y15-24","PL62",1999,45.2,"Warminsko-Mazurskie"
"Y15-24","PL63",1999,16.4,"Pomorskie"
"Y15-24","PT",1999,9.1,"Portugal"
"Y15-24","PT1",1999,9.3,"Continente"
"Y15-24","PT11",1999,7.7,"Norte"
"Y15-24","PT15",1999,NA,"Algarve"
"Y15-24","PT16",1999,6.5,"Centro (PT)"
"Y15-24","PT17",1999,12.9,"Área Metropolitana de Lisboa"
"Y15-24","PT18",1999,NA,"Alentejo"
"Y15-24","PT2",1999,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT20",1999,NA,"Região Autónoma dos Açores (PT)"
"Y15-24","PT3",1999,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","PT30",1999,NA,"Região Autónoma da Madeira (PT)"
"Y15-24","RO",1999,17.3,"Romania"
"Y15-24","RO1",1999,18.7,"Macroregiunea unu"
"Y15-24","RO11",1999,18.6,"Nord-Vest"
"Y15-24","RO12",1999,18.8,"Centru"
"Y15-24","RO2",1999,16.8,"Macroregiunea doi"
"Y15-24","RO21",1999,16.5,"Nord-Est"
"Y15-24","RO22",1999,17.1,"Sud-Est"
"Y15-24","RO3",1999,20.4,"Macroregiunea trei"
"Y15-24","RO31",1999,20,"Sud - Muntenia"
"Y15-24","RO32",1999,21.3,"Bucuresti - Ilfov"
"Y15-24","RO4",1999,12.5,"Macroregiunea patru"
"Y15-24","RO41",1999,11.4,"Sud-Vest Oltenia"
"Y15-24","RO42",1999,13.7,"Vest"
"Y15-24","SE",1999,16.3,"Sweden"
"Y15-24","SE1",1999,14.9,"Östra Sverige"
"Y15-24","SE11",1999,NA,"Stockholm"
"Y15-24","SE12",1999,20.9,"Östra Mellansverige"
"Y15-24","SE2",1999,16.3,"Södra Sverige"
"Y15-24","SE21",1999,NA,"Småland med öarna"
"Y15-24","SE22",1999,20.5,"Sydsverige"
"Y15-24","SE23",1999,14.7,"Västsverige"
"Y15-24","SE3",1999,19.1,"Norra Sverige"
"Y15-24","SE31",1999,23.5,"Norra Mellansverige"
"Y15-24","SE32",1999,NA,"Mellersta Norrland"
"Y15-24","SE33",1999,NA,"Övre Norrland"
"Y15-24","SI",1999,18.5,"Slovenia"
"Y15-24","SI0",1999,18.5,"Slovenija"
"Y15-24","SK",1999,32,"Slovakia"
"Y15-24","SK0",1999,32,"Slovensko"
"Y15-24","SK01",1999,16.7,"Bratislavský kraj"
"Y15-24","SK02",1999,27.9,"Západné Slovensko"
"Y15-24","SK03",1999,35.7,"Stredné Slovensko"
"Y15-24","SK04",1999,39,"Východné Slovensko"
"Y15-24","UK",1999,12.4,"United Kingdom"
"Y15-24","UKC",1999,18.4,"North East (UK)"
"Y15-24","UKC1",1999,19.6,"Tees Valley and Durham"
"Y15-24","UKC2",1999,17.4,"Northumberland and Tyne and Wear"
"Y15-24","UKD",1999,13.7,"North West (UK)"
"Y15-24","UKD1",1999,NA,"Cumbria"
"Y15-24","UKD3",1999,15.7,"Greater Manchester"
"Y15-24","UKD4",1999,NA,"Lancashire"
"Y15-24","UKE",1999,12,"Yorkshire and The Humber"
"Y15-24","UKE1",1999,18.8,"East Yorkshire and Northern Lincolnshire"
"Y15-24","UKE2",1999,NA,"North Yorkshire"
"Y15-24","UKE3",1999,14,"South Yorkshire"
"Y15-24","UKE4",1999,9.6,"West Yorkshire"
"Y15-24","UKF",1999,13.7,"East Midlands (UK)"
"Y15-24","UKF1",1999,14.2,"Derbyshire and Nottinghamshire"
"Y15-24","UKF2",1999,13,"Leicestershire, Rutland and Northamptonshire"
"Y15-24","UKF3",1999,NA,"Lincolnshire"
"Y15-24","UKG",1999,13.7,"West Midlands (UK)"
"Y15-24","UKG1",1999,NA,"Herefordshire, Worcestershire and Warwickshire"
"Y15-24","UKG2",1999,13.4,"Shropshire and Staffordshire"
"Y15-24","UKG3",1999,14.9,"West Midlands"
"Y15-24","UKH",1999,8.7,"East of England"
"Y15-24","UKH1",1999,8.5,"East Anglia"
"Y15-24","UKH2",1999,11.2,"Bedfordshire and Hertfordshire"
"Y15-24","UKH3",1999,NA,"Essex"
"Y15-24","UKI",1999,13.7,"London"
"Y15-24","UKI1",1999,16.3,"Inner London (NUTS 2010)"
"Y15-24","UKI2",1999,12.1,"Outer London (NUTS 2010)"
"Y15-24","UKJ",1999,7,"South East (UK)"
"Y15-24","UKJ1",1999,NA,"Berkshire, Buckinghamshire and Oxfordshire"
"Y15-24","UKJ2",1999,6.1,"Surrey, East and West Sussex"
"Y15-24","UKJ3",1999,11.4,"Hampshire and Isle of Wight"
"Y15-24","UKJ4",1999,10.3,"Kent"
"Y15-24","UKK",1999,11.1,"South West (UK)"
"Y15-24","UKK1",1999,8.2,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y15-24","UKK2",1999,NA,"Dorset and Somerset"
"Y15-24","UKK3",1999,NA,"Cornwall and Isles of Scilly"
"Y15-24","UKK4",1999,15.3,"Devon"
"Y15-24","UKL",1999,16.8,"Wales"
"Y15-24","UKL1",1999,16.4,"West Wales and The Valleys"
"Y15-24","UKL2",1999,17.5,"East Wales"
"Y15-24","UKM",1999,16,"Scotland"
"Y15-24","UKM2",1999,16.7,"Eastern Scotland"
"Y15-24","UKM3",1999,18.5,"South Western Scotland"
"Y15-24","UKN",1999,10.3,"Northern Ireland (UK)"
"Y15-24","UKN0",1999,10.3,"Northern Ireland (UK)"
"Y20-64","AT",1999,4.6,"Austria"
"Y20-64","AT1",1999,5.4,"Ostösterreich"
"Y20-64","AT11",1999,4.8,"Burgenland (AT)"
"Y20-64","AT12",1999,4.2,"Niederösterreich"
"Y20-64","AT13",1999,6.5,"Wien"
"Y20-64","AT2",1999,4.1,"Südösterreich"
"Y20-64","AT21",1999,4.1,"Kärnten"
"Y20-64","AT22",1999,4.1,"Steiermark"
"Y20-64","AT3",1999,4,"Westösterreich"
"Y20-64","AT31",1999,4.7,"Oberösterreich"
"Y20-64","AT32",1999,3,"Salzburg"
"Y20-64","AT33",1999,3.3,"Tirol"
"Y20-64","AT34",1999,4.2,"Vorarlberg"
"Y20-64","BE",1999,8.4,"Belgium"
"Y20-64","BE1",1999,15.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE10",1999,15.6,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y20-64","BE2",1999,5.4,"Vlaams Gewest"
"Y20-64","BE21",1999,6.3,"Prov. Antwerpen"
"Y20-64","BE22",1999,6.3,"Prov. Limburg (BE)"
"Y20-64","BE23",1999,6.3,"Prov. Oost-Vlaanderen"
"Y20-64","BE24",1999,3.5,"Prov. Vlaams-Brabant"
"Y20-64","BE25",1999,3.9,"Prov. West-Vlaanderen"
"Y20-64","BE3",1999,12.2,"Région wallonne"
"Y20-64","BE31",1999,7.6,"Prov. Brabant Wallon"
"Y20-64","BE32",1999,15.9,"Prov. Hainaut"
"Y20-64","BE33",1999,11.9,"Prov. Liège"
"Y20-64","BE34",1999,6.7,"Prov. Luxembourg (BE)"
"Y20-64","BE35",1999,9.7,"Prov. Namur"
"Y20-64","CH",1999,2.9,"Switzerland"
"Y20-64","CH0",1999,2.9,"Schweiz/Suisse/Svizzera"
"Y20-64","CZ",1999,7.9,"Czech Republic"
"Y20-64","CZ0",1999,7.9,"Ceská republika"
"Y20-64","CZ01",1999,3.3,"Praha"
"Y20-64","CZ02",1999,7.3,"Strední Cechy"
"Y20-64","CZ03",1999,5.9,"Jihozápad"
"Y20-64","CZ04",1999,12.2,"Severozápad"
"Y20-64","CZ05",1999,7.1,"Severovýchod"
"Y20-64","CZ06",1999,7.3,"Jihovýchod"
"Y20-64","CZ07",1999,9,"Strední Morava"
"Y20-64","CZ08",1999,11.8,"Moravskoslezsko"
"Y20-64","DE",1999,9,"Germany (until 1990 former territory of the FRG)"
"Y20-64","DE1",1999,5.5,"Baden-Württemberg"
"Y20-64","DE11",1999,5.4,"Stuttgart"
"Y20-64","DE12",1999,6.3,"Karlsruhe"
"Y20-64","DE13",1999,5.4,"Freiburg"
"Y20-64","DE14",1999,4.7,"Tübingen"
"Y20-64","DE2",1999,5,"Bayern"
"Y20-64","DE21",1999,4.1,"Oberbayern"
"Y20-64","DE22",1999,5,"Niederbayern"
"Y20-64","DE23",1999,4.6,"Oberpfalz"
"Y20-64","DE24",1999,6.3,"Oberfranken"
"Y20-64","DE25",1999,6.5,"Mittelfranken"
"Y20-64","DE26",1999,6,"Unterfranken"
"Y20-64","DE27",1999,4.7,"Schwaben"
"Y20-64","DE3",1999,15.2,"Berlin"
"Y20-64","DE30",1999,15.2,"Berlin"
"Y20-64","DE4",1999,16.2,"Brandenburg"
"Y20-64","DE40",1999,16.2,"Brandenburg"
"Y20-64","DE5",1999,11.7,"Bremen"
"Y20-64","DE50",1999,11.7,"Bremen"
"Y20-64","DE6",1999,8.7,"Hamburg"
"Y20-64","DE60",1999,8.7,"Hamburg"
"Y20-64","DE7",1999,7.3,"Hessen"
"Y20-64","DE71",1999,6.9,"Darmstadt"
"Y20-64","DE72",1999,7.5,"Gießen"
"Y20-64","DE73",1999,8.6,"Kassel"
"Y20-64","DE8",1999,19.1,"Mecklenburg-Vorpommern"
"Y20-64","DE80",1999,19.1,"Mecklenburg-Vorpommern"
"Y20-64","DE9",1999,7.4,"Niedersachsen"
"Y20-64","DE91",1999,8.9,"Braunschweig"
"Y20-64","DE92",1999,8.1,"Hannover"
"Y20-64","DE93",1999,6.6,"Lüneburg"
"Y20-64","DE94",1999,6.4,"Weser-Ems"
"Y20-64","DEA",1999,7.5,"Nordrhein-Westfalen"
"Y20-64","DEA1",1999,7.7,"Düsseldorf"
"Y20-64","DEA2",1999,6.8,"Köln"
"Y20-64","DEA3",1999,7.5,"Münster"
"Y20-64","DEA4",1999,6.5,"Detmold"
"Y20-64","DEA5",1999,8.4,"Arnsberg"
"Y20-64","DEB",1999,6.1,"Rheinland-Pfalz"
"Y20-64","DEB1",1999,6,"Koblenz"
"Y20-64","DEB2",1999,6,"Trier"
"Y20-64","DEB3",1999,6.3,"Rheinhessen-Pfalz"
"Y20-64","DEC",1999,7.5,"Saarland"
"Y20-64","DEC0",1999,7.5,"Saarland"
"Y20-64","DED",1999,16.7,"Sachsen"
"Y20-64","DEE",1999,21.6,"Sachsen-Anhalt"
"Y20-64","DEE0",1999,21.6,"Sachsen-Anhalt"
"Y20-64","DEF",1999,7.6,"Schleswig-Holstein"
"Y20-64","DEF0",1999,7.6,"Schleswig-Holstein"
"Y20-64","DEG",1999,15.1,"Thüringen"
"Y20-64","DEG0",1999,15.1,"Thüringen"
"Y20-64","DK",1999,4.9,"Denmark"
"Y20-64","DK0",1999,4.9,"Danmark"
"Y20-64","EE",1999,11.2,"Estonia"
"Y20-64","EE0",1999,11.2,"Eesti"
"Y20-64","EE00",1999,11.2,"Eesti"
"Y20-64","EL",1999,11.3,"Greece"
"Y20-64","EL1",1999,12,"Voreia Ellada (NUTS 2010)"
"Y20-64","EL11",1999,12.5,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y20-64","EL12",1999,11.4,"Kentriki Makedonia (NUTS 2010)"
"Y20-64","EL13",1999,13.2,"Dytiki Makedonia (NUTS 2010)"
"Y20-64","EL14",1999,12.6,"Thessalia (NUTS 2010)"
"Y20-64","EL2",1999,11,"Kentriki Ellada (NUTS 2010)"
"Y20-64","EL21",1999,14,"Ipeiros (NUTS 2010)"
"Y20-64","EL22",1999,5.9,"Ionia Nisia (NUTS 2010)"
"Y20-64","EL23",1999,11.3,"Dytiki Ellada (NUTS 2010)"
"Y20-64","EL24",1999,14.5,"Sterea Ellada (NUTS 2010)"
"Y20-64","EL25",1999,7.5,"Peloponnisos (NUTS 2010)"
"Y20-64","EL3",1999,11.9,"Attiki"
"Y20-64","EL30",1999,11.9,"Attiki"
"Y20-64","EL4",1999,8,"Nisia Aigaiou, Kriti"
"Y20-64","EL41",1999,11.4,"Voreio Aigaio"
"Y20-64","EL42",1999,7.3,"Notio Aigaio"
"Y20-64","EL43",1999,7.4,"Kriti"
"Y20-64","ES",1999,14.8,"Spain"
"Y20-64","ES1",1999,16.1,"Noroeste (ES)"
"Y20-64","ES11",1999,16,"Galicia"
"Y20-64","ES12",1999,17.3,"Principado de Asturias"
"Y20-64","ES13",1999,14.8,"Cantabria"
"Y20-64","ES2",1999,11.3,"Noreste (ES)"
"Y20-64","ES21",1999,13.6,"País Vasco"
"Y20-64","ES22",1999,8.1,"Comunidad Foral de Navarra"
"Y20-64","ES23",1999,6.3,"La Rioja"
"Y20-64","ES24",1999,9.6,"Aragón"
"Y20-64","ES3",1999,12.3,"Comunidad de Madrid"
"Y20-64","ES30",1999,12.3,"Comunidad de Madrid"
"Y20-64","ES4",1999,16.5,"Centro (ES)"
"Y20-64","ES41",1999,14.7,"Castilla y León"
"Y20-64","ES42",1999,14.6,"Castilla-la Mancha"
"Y20-64","ES43",1999,24.1,"Extremadura"
"Y20-64","ES5",1999,10.7,"Este (ES)"
"Y20-64","ES51",1999,9.9,"Cataluña"
"Y20-64","ES52",1999,12.9,"Comunidad Valenciana"
"Y20-64","ES53",1999,6.8,"Illes Balears"
"Y20-64","ES6",1999,23.2,"Sur (ES)"
"Y20-64","ES61",1999,24.9,"Andalucía"
"Y20-64","ES62",1999,13.2,"Región de Murcia"
"Y20-64","ES63",1999,23.9,"Ciudad Autónoma de Ceuta (ES)"
"Y20-64","ES64",1999,20.7,"Ciudad Autónoma de Melilla (ES)"
"Y20-64","ES7",1999,12.9,"Canarias (ES)"
"Y20-64","ES70",1999,12.9,"Canarias (ES)"
"Y20-64","EU15",1999,9.1,"European Union (15 countries)"
"Y20-64","FI",1999,9.8,"Finland"
"Y20-64","FI1",1999,9.9,"Manner-Suomi"
"Y20-64","FI19",1999,10.6,"Länsi-Suomi"
"Y20-64","FI2",1999,NA,"Åland"
"Y20-64","FI20",1999,NA,"Åland"
"Y20-64","FR",1999,11.6,"France"
"Y20-64","FR1",1999,10.2,"Île de France"
"Y20-64","FR10",1999,10.2,"Île de France"
"Y20-64","FR2",1999,11.5,"Bassin Parisien"
"Y20-64","FR21",1999,12.5,"Champagne-Ardenne"
"Y20-64","FR22",1999,12.9,"Picardie"
"Y20-64","FR23",1999,13.6,"Haute-Normandie"
"Y20-64","FR24",1999,10.5,"Centre (FR)"
"Y20-64","FR25",1999,9.5,"Basse-Normandie"
"Y20-64","FR26",1999,10.1,"Bourgogne"
"Y20-64","FR3",1999,17.3,"Nord - Pas-de-Calais"
"Y20-64","FR30",1999,17.3,"Nord - Pas-de-Calais"
"Y20-64","FR4",1999,9.3,"Est (FR)"
"Y20-64","FR41",1999,10.9,"Lorraine"
"Y20-64","FR42",1999,7.2,"Alsace"
"Y20-64","FR43",1999,9.6,"Franche-Comté"
"Y20-64","FR5",1999,10.6,"Ouest (FR)"
"Y20-64","FR51",1999,11.9,"Pays de la Loire"
"Y20-64","FR52",1999,9.3,"Bretagne"
"Y20-64","FR53",1999,10.3,"Poitou-Charentes"
"Y20-64","FR6",1999,11.1,"Sud-Ouest (FR)"
"Y20-64","FR61",1999,11.6,"Aquitaine"
"Y20-64","FR62",1999,10.9,"Midi-Pyrénées"
"Y20-64","FR63",1999,9.4,"Limousin"
"Y20-64","FR7",1999,9.7,"Centre-Est (FR)"
"Y20-64","FR71",1999,9.6,"Rhône-Alpes"
"Y20-64","FR72",1999,10.4,"Auvergne"
"Y20-64","FR8",1999,17.1,"Méditerranée"
"Y20-64","FR81",1999,16.9,"Languedoc-Roussillon"
"Y20-64","FR82",1999,16.7,"Provence-Alpes-Côte d'Azur"
"Y20-64","FR83",1999,25.1,"Corse"
"Y20-64","HU",1999,6.6,"Hungary"
"Y20-64","HU1",1999,4.7,"Közép-Magyarország"
"Y20-64","HU10",1999,4.7,"Közép-Magyarország"
"Y20-64","HU2",1999,6,"Dunántúl"
"Y20-64","HU21",1999,5.8,"Közép-Dunántúl"
"Y20-64","HU22",1999,4.3,"Nyugat-Dunántúl"
"Y20-64","HU23",1999,8,"Dél-Dunántúl"
"Y20-64","HU3",1999,8.7,"Alföld és Észak"
"Y20-64","HU31",1999,11,"Észak-Magyarország"
"Y20-64","HU32",1999,9.8,"Észak-Alföld"
"Y20-64","HU33",1999,5.5,"Dél-Alföld"
"Y20-64","IE",1999,5.6,"Ireland"
"Y20-64","IE0",1999,5.6,"Éire/Ireland"
"Y20-64","IE01",1999,6.7,"Border, Midland and Western"
"Y20-64","IE02",1999,5.2,"Southern and Eastern"
"Y20-64","IS",1999,2,"Iceland"
"Y20-64","IS0",1999,2,"Ísland"
"Y20-64","IS00",1999,2,"Ísland"
"Y20-64","IT",1999,11.2,"Italy"
"Y20-64","ITC",1999,5.9,"Nord-Ovest"
"Y20-64","ITC1",1999,7.3,"Piemonte"
"Y20-64","ITC2",1999,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y20-64","ITC3",1999,10.3,"Liguria"
"Y20-64","ITC4",1999,4.5,"Lombardia"
"Y20-64","ITF",1999,20.2,"Sud"
"Y20-64","ITF1",1999,10.1,"Abruzzo"
"Y20-64","ITF2",1999,15.4,"Molise"
"Y20-64","ITF3",1999,22.1,"Campania"
"Y20-64","ITF4",1999,18.4,"Puglia"
"Y20-64","ITF5",1999,16.2,"Basilicata"
"Y20-64","ITF6",1999,27.2,"Calabria"
"Y20-64","ITG",1999,22.4,"Isole"
"Y20-64","ITG1",1999,23,"Sicilia"
"Y20-64","ITG2",1999,20.5,"Sardegna"
"Y20-64","ITH",1999,4.6,"Nord-Est"
"Y20-64","ITH1",1999,2.2,"Provincia Autonoma di Bolzano/Bozen"
"Y20-64","ITH2",1999,5.2,"Provincia Autonoma di Trento"
"Y20-64","ITH3",1999,4.7,"Veneto"
"Y20-64","ITH4",1999,5.1,"Friuli-Venezia Giulia"
"Y20-64","ITI",1999,9.8,"Centro (IT)"
"Y20-64","ITI1",1999,7.9,"Toscana"
"Y20-64","ITI2",1999,6.8,"Umbria"
"Y20-64","ITI4",1999,12.7,"Lazio"
"Y20-64","LT",1999,13.1,"Lithuania"
"Y20-64","LT0",1999,13.1,"Lietuva"
"Y20-64","LT00",1999,13.1,"Lietuva"
"Y20-64","LU",1999,2.2,"Luxembourg"
"Y20-64","LU0",1999,2.2,"Luxembourg"
"Y20-64","LU00",1999,2.2,"Luxembourg"
"Y20-64","LV",1999,13.5,"Latvia"
"Y20-64","LV0",1999,13.5,"Latvija"
"Y20-64","LV00",1999,13.5,"Latvija"
"Y20-64","NL",1999,3.1,"Netherlands"
"Y20-64","NL1",1999,5.2,"Noord-Nederland"
"Y20-64","NL11",1999,5.3,"Groningen"
"Y20-64","NL12",1999,3.4,"Friesland (NL)"
"Y20-64","NL13",1999,7.4,"Drenthe"
"Y20-64","NL2",1999,2.7,"Oost-Nederland"
"Y20-64","NL21",1999,2.4,"Overijssel"
"Y20-64","NL22",1999,2.7,"Gelderland"
"Y20-64","NL23",1999,3.9,"Flevoland"
"Y20-64","NL3",1999,3,"West-Nederland"
"Y20-64","NL31",1999,2.7,"Utrecht"
"Y20-64","NL32",1999,3.2,"Noord-Holland"
"Y20-64","NL33",1999,2.8,"Zuid-Holland"
"Y20-64","NL34",1999,5.2,"Zeeland"
"Y20-64","NL4",1999,2.5,"Zuid-Nederland"
"Y20-64","NL41",1999,2.3,"Noord-Brabant"
"Y20-64","NL42",1999,2.9,"Limburg (NL)"
"Y20-64","NO",1999,2.4,"Norway"
"Y20-64","NO0",1999,2.4,"Norge"
"Y20-64","NO01",1999,1.7,"Oslo og Akershus"
"Y20-64","NO02",1999,2.3,"Hedmark og Oppland"
"Y20-64","NO03",1999,2.8,"Sør-Østlandet"
"Y20-64","NO04",1999,2.5,"Agder og Rogaland"
"Y20-64","NO05",1999,2.1,"Vestlandet"
"Y20-64","NO06",1999,2.8,"Trøndelag"
"Y20-64","NO07",1999,3.2,"Nord-Norge"
"Y20-64","PL",1999,12.3,"Poland"
"Y20-64","PL1",1999,11,"Region Centralny"
"Y20-64","PL11",1999,12.4,"Lódzkie"
"Y20-64","PL12",1999,10.2,"Mazowieckie"
"Y20-64","PL2",1999,10.2,"Region Poludniowy"
"Y20-64","PL21",1999,9.4,"Malopolskie"
"Y20-64","PL22",1999,10.9,"Slaskie"
"Y20-64","PL3",1999,12.5,"Region Wschodni"
"Y20-64","PL31",1999,11.3,"Lubelskie"
"Y20-64","PL32",1999,12.7,"Podkarpackie"
"Y20-64","PL33",1999,13.9,"Swietokrzyskie"
"Y20-64","PL34",1999,12.6,"Podlaskie"
"Y20-64","PL4",1999,13.4,"Region Pólnocno-Zachodni"
"Y20-64","PL41",1999,9.5,"Wielkopolskie"
"Y20-64","PL42",1999,19.3,"Zachodniopomorskie"
"Y20-64","PL43",1999,15.8,"Lubuskie"
"Y20-64","PL5",1999,14.5,"Region Poludniowo-Zachodni"
"Y20-64","PL51",1999,14.8,"Dolnoslaskie"
"Y20-64","PL52",1999,13.7,"Opolskie"
"Y20-64","PL6",1999,13.9,"Region Pólnocny"
"Y20-64","PL61",1999,13.1,"Kujawsko-Pomorskie"
"Y20-64","PL62",1999,19.3,"Warminsko-Mazurskie"
"Y20-64","PL63",1999,11.1,"Pomorskie"
"Y20-64","PT",1999,4.7,"Portugal"
"Y20-64","PT1",1999,4.8,"Continente"
"Y20-64","PT11",1999,4.6,"Norte"
"Y20-64","PT15",1999,NA,"Algarve"
"Y20-64","PT16",1999,2.6,"Centro (PT)"
"Y20-64","PT17",1999,6.2,"Área Metropolitana de Lisboa"
"Y20-64","PT18",1999,7.4,"Alentejo"
"Y20-64","PT2",1999,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT20",1999,NA,"Região Autónoma dos Açores (PT)"
"Y20-64","PT3",1999,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","PT30",1999,NA,"Região Autónoma da Madeira (PT)"
"Y20-64","RO",1999,6.2,"Romania"
"Y20-64","RO1",1999,6.5,"Macroregiunea unu"
"Y20-64","RO11",1999,6.5,"Nord-Vest"
"Y20-64","RO12",1999,6.5,"Centru"
"Y20-64","RO2",1999,7.2,"Macroregiunea doi"
"Y20-64","RO21",1999,7.3,"Nord-Est"
"Y20-64","RO22",1999,7,"Sud-Est"
"Y20-64","RO3",1999,5.6,"Macroregiunea trei"
"Y20-64","RO31",1999,6.4,"Sud - Muntenia"
"Y20-64","RO32",1999,4.5,"Bucuresti - Ilfov"
"Y20-64","RO4",1999,5.4,"Macroregiunea patru"
"Y20-64","RO41",1999,4.4,"Sud-Vest Oltenia"
"Y20-64","RO42",1999,6.6,"Vest"
"Y20-64","SE",1999,7.4,"Sweden"
"Y20-64","SE1",1999,5.6,"Östra Sverige"
"Y20-64","SE11",1999,3.7,"Stockholm"
"Y20-64","SE12",1999,7.9,"Östra Mellansverige"
"Y20-64","SE2",1999,7.4,"Södra Sverige"
"Y20-64","SE21",1999,7.1,"Småland med öarna"
"Y20-64","SE22",1999,8.4,"Sydsverige"
"Y20-64","SE23",1999,6.8,"Västsverige"
"Y20-64","SE3",1999,10.6,"Norra Sverige"
"Y20-64","SE31",1999,11.3,"Norra Mellansverige"
"Y20-64","SE32",1999,8,"Mellersta Norrland"
"Y20-64","SE33",1999,11.5,"Övre Norrland"
"Y20-64","SI",1999,7.1,"Slovenia"
"Y20-64","SI0",1999,7.1,"Slovenija"
"Y20-64","SK",1999,14.5,"Slovakia"
"Y20-64","SK0",1999,14.5,"Slovensko"
"Y20-64","SK01",1999,6.3,"Bratislavský kraj"
"Y20-64","SK02",1999,12.8,"Západné Slovensko"
"Y20-64","SK03",1999,16.4,"Stredné Slovensko"
"Y20-64","SK04",1999,18.7,"Východné Slovensko"
"Y20-64","UK",1999,5.5,"United Kingdom"
"Y20-64","UKC",1999,9.5,"North East (UK)"
"Y20-64","UKC1",1999,9.7,"Tees Valley and Durham"
"Y20-64","UKC2",1999,9.3,"Northumberland and Tyne and Wear"
"Y20-64","UKD",1999,5.5,"North West (UK)"
"Y20-64","UKD1",1999,6.1,"Cumbria"
"Y20-64","UKD3",1999,5.6,"Greater Manchester"
"Y20-64","UKD4",1999,3.7,"Lancashire"
"Y20-64","UKE",1999,6,"Yorkshire and The Humber"
"Y20-64","UKE1",1999,7.5,"East Yorkshire and Northern Lincolnshire"
"Y20-64","UKE2",1999,3.2,"North Yorkshire"
"Y20-64","UKE3",1999,7,"South Yorkshire"
"Y20-64","UKE4",1999,5.6,"West Yorkshire"
"Y20-64","UKF",1999,4.4,"East Midlands (UK)"
"Y20-64","UKF1",1999,4.9,"Derbyshire and Nottinghamshire"
"Y20-64","UKF2",1999,3.9,"Leicestershire, Rutland and Northamptonshire"
"Y20-64","UKF3",1999,3.8,"Lincolnshire"
"Y20-64","UKG",1999,6.1,"West Midlands (UK)"
"Y20-64","UKG1",1999,4.4,"Herefordshire, Worcestershire and Warwickshire"
"Y20-64","UKG2",1999,5.4,"Shropshire and Staffordshire"
"Y20-64","UKG3",1999,7.4,"West Midlands"
"Y20-64","UKH",1999,3.9,"East of England"
"Y20-64","UKH1",1999,3.8,"East Anglia"
"Y20-64","UKH2",1999,3.9,"Bedfordshire and Hertfordshire"
"Y20-64","UKH3",1999,3.9,"Essex"
"Y20-64","UKI",1999,7.1,"London"
"Y20-64","UKI1",1999,8.7,"Inner London (NUTS 2010)"
"Y20-64","UKI2",1999,6.2,"Outer London (NUTS 2010)"
"Y20-64","UKJ",1999,3.3,"South East (UK)"
"Y20-64","UKJ1",1999,2.5,"Berkshire, Buckinghamshire and Oxfordshire"
"Y20-64","UKJ2",1999,3.3,"Surrey, East and West Sussex"
"Y20-64","UKJ3",1999,4,"Hampshire and Isle of Wight"
"Y20-64","UKJ4",1999,3.6,"Kent"
"Y20-64","UKK",1999,4.3,"South West (UK)"
"Y20-64","UKK1",1999,3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y20-64","UKK2",1999,4.4,"Dorset and Somerset"
"Y20-64","UKK3",1999,7.3,"Cornwall and Isles of Scilly"
"Y20-64","UKK4",1999,5.8,"Devon"
"Y20-64","UKL",1999,6.1,"Wales"
"Y20-64","UKL1",1999,6.8,"West Wales and The Valleys"
"Y20-64","UKL2",1999,5.2,"East Wales"
"Y20-64","UKM",1999,6.7,"Scotland"
"Y20-64","UKM2",1999,6,"Eastern Scotland"
"Y20-64","UKM3",1999,7.8,"South Western Scotland"
"Y20-64","UKN",1999,6.9,"Northern Ireland (UK)"
"Y20-64","UKN0",1999,6.9,"Northern Ireland (UK)"
"Y_GE15","AT",1999,4.7,"Austria"
"Y_GE15","AT1",1999,5.5,"Ostösterreich"
"Y_GE15","AT11",1999,4.9,"Burgenland (AT)"
"Y_GE15","AT12",1999,4.3,"Niederösterreich"
"Y_GE15","AT13",1999,6.7,"Wien"
"Y_GE15","AT2",1999,4.2,"Südösterreich"
"Y_GE15","AT21",1999,4,"Kärnten"
"Y_GE15","AT22",1999,4.2,"Steiermark"
"Y_GE15","AT3",1999,4,"Westösterreich"
"Y_GE15","AT31",1999,4.7,"Oberösterreich"
"Y_GE15","AT32",1999,3.1,"Salzburg"
"Y_GE15","AT33",1999,3.3,"Tirol"
"Y_GE15","AT34",1999,4.5,"Vorarlberg"
"Y_GE15","BE",1999,8.6,"Belgium"
"Y_GE15","BE1",1999,15.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE10",1999,15.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE15","BE2",1999,5.6,"Vlaams Gewest"
"Y_GE15","BE21",1999,6.5,"Prov. Antwerpen"
"Y_GE15","BE22",1999,6.6,"Prov. Limburg (BE)"
"Y_GE15","BE23",1999,6.6,"Prov. Oost-Vlaanderen"
"Y_GE15","BE24",1999,3.7,"Prov. Vlaams-Brabant"
"Y_GE15","BE25",1999,4.1,"Prov. West-Vlaanderen"
"Y_GE15","BE3",1999,12.3,"Région wallonne"
"Y_GE15","BE31",1999,8,"Prov. Brabant Wallon"
"Y_GE15","BE32",1999,16,"Prov. Hainaut"
"Y_GE15","BE33",1999,12,"Prov. Liège"
"Y_GE15","BE34",1999,6.8,"Prov. Luxembourg (BE)"
"Y_GE15","BE35",1999,10,"Prov. Namur"
"Y_GE15","CH",1999,3.1,"Switzerland"
"Y_GE15","CH0",1999,3.1,"Schweiz/Suisse/Svizzera"
"Y_GE15","CZ",1999,8.5,"Czech Republic"
"Y_GE15","CZ0",1999,8.5,"Ceská republika"
"Y_GE15","CZ01",1999,3.6,"Praha"
"Y_GE15","CZ02",1999,8,"Strední Cechy"
"Y_GE15","CZ03",1999,6.2,"Jihozápad"
"Y_GE15","CZ04",1999,13.1,"Severozápad"
"Y_GE15","CZ05",1999,7.6,"Severovýchod"
"Y_GE15","CZ06",1999,8,"Jihovýchod"
"Y_GE15","CZ07",1999,9.6,"Strední Morava"
"Y_GE15","CZ08",1999,12.5,"Moravskoslezsko"
"Y_GE15","DE",1999,8.9,"Germany (until 1990 former territory of the FRG)"
"Y_GE15","DE1",1999,5.4,"Baden-Württemberg"
"Y_GE15","DE11",1999,5.3,"Stuttgart"
"Y_GE15","DE12",1999,6.2,"Karlsruhe"
"Y_GE15","DE13",1999,5.3,"Freiburg"
"Y_GE15","DE14",1999,4.7,"Tübingen"
"Y_GE15","DE2",1999,5,"Bayern"
"Y_GE15","DE21",1999,4,"Oberbayern"
"Y_GE15","DE22",1999,4.9,"Niederbayern"
"Y_GE15","DE23",1999,4.6,"Oberpfalz"
"Y_GE15","DE24",1999,6.3,"Oberfranken"
"Y_GE15","DE25",1999,6.6,"Mittelfranken"
"Y_GE15","DE26",1999,6.3,"Unterfranken"
"Y_GE15","DE27",1999,4.6,"Schwaben"
"Y_GE15","DE3",1999,15.3,"Berlin"
"Y_GE15","DE30",1999,15.3,"Berlin"
"Y_GE15","DE4",1999,15.8,"Brandenburg"
"Y_GE15","DE40",1999,15.8,"Brandenburg"
"Y_GE15","DE5",1999,11.5,"Bremen"
"Y_GE15","DE50",1999,11.5,"Bremen"
"Y_GE15","DE6",1999,8.6,"Hamburg"
"Y_GE15","DE60",1999,8.6,"Hamburg"
"Y_GE15","DE7",1999,7.3,"Hessen"
"Y_GE15","DE71",1999,6.9,"Darmstadt"
"Y_GE15","DE72",1999,7.5,"Gießen"
"Y_GE15","DE73",1999,8.4,"Kassel"
"Y_GE15","DE8",1999,18.2,"Mecklenburg-Vorpommern"
"Y_GE15","DE80",1999,18.2,"Mecklenburg-Vorpommern"
"Y_GE15","DE9",1999,7.4,"Niedersachsen"
"Y_GE15","DE91",1999,8.8,"Braunschweig"
"Y_GE15","DE92",1999,8,"Hannover"
"Y_GE15","DE93",1999,6.4,"Lüneburg"
"Y_GE15","DE94",1999,6.4,"Weser-Ems"
"Y_GE15","DEA",1999,7.5,"Nordrhein-Westfalen"
"Y_GE15","DEA1",1999,7.7,"Düsseldorf"
"Y_GE15","DEA2",1999,6.8,"Köln"
"Y_GE15","DEA3",1999,7.6,"Münster"
"Y_GE15","DEA4",1999,6.4,"Detmold"
"Y_GE15","DEA5",1999,8.3,"Arnsberg"
"Y_GE15","DEB",1999,6.1,"Rheinland-Pfalz"
"Y_GE15","DEB1",1999,6,"Koblenz"
"Y_GE15","DEB2",1999,5.7,"Trier"
"Y_GE15","DEB3",1999,6.2,"Rheinhessen-Pfalz"
"Y_GE15","DEC",1999,7.2,"Saarland"
"Y_GE15","DEC0",1999,7.2,"Saarland"
"Y_GE15","DED",1999,16,"Sachsen"
"Y_GE15","DEE",1999,20.8,"Sachsen-Anhalt"
"Y_GE15","DEE0",1999,20.8,"Sachsen-Anhalt"
"Y_GE15","DEF",1999,7.7,"Schleswig-Holstein"
"Y_GE15","DEF0",1999,7.7,"Schleswig-Holstein"
"Y_GE15","DEG",1999,14.5,"Thüringen"
"Y_GE15","DEG0",1999,14.5,"Thüringen"
"Y_GE15","DK",1999,5.1,"Denmark"
"Y_GE15","DK0",1999,5.1,"Danmark"
"Y_GE15","EE",1999,11.6,"Estonia"
"Y_GE15","EE0",1999,11.6,"Eesti"
"Y_GE15","EE00",1999,11.6,"Eesti"
"Y_GE15","EL",1999,11.9,"Greece"
"Y_GE15","EL1",1999,12.5,"Voreia Ellada (NUTS 2010)"
"Y_GE15","EL11",1999,13,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE15","EL12",1999,11.8,"Kentriki Makedonia (NUTS 2010)"
"Y_GE15","EL13",1999,14.4,"Dytiki Makedonia (NUTS 2010)"
"Y_GE15","EL14",1999,13.1,"Thessalia (NUTS 2010)"
"Y_GE15","EL2",1999,11.5,"Kentriki Ellada (NUTS 2010)"
"Y_GE15","EL21",1999,14.2,"Ipeiros (NUTS 2010)"
"Y_GE15","EL22",1999,5.8,"Ionia Nisia (NUTS 2010)"
"Y_GE15","EL23",1999,12,"Dytiki Ellada (NUTS 2010)"
"Y_GE15","EL24",1999,15.2,"Sterea Ellada (NUTS 2010)"
"Y_GE15","EL25",1999,7.9,"Peloponnisos (NUTS 2010)"
"Y_GE15","EL3",1999,12.6,"Attiki"
"Y_GE15","EL30",1999,12.6,"Attiki"
"Y_GE15","EL4",1999,8.2,"Nisia Aigaiou, Kriti"
"Y_GE15","EL41",1999,11.7,"Voreio Aigaio"
"Y_GE15","EL42",1999,7.6,"Notio Aigaio"
"Y_GE15","EL43",1999,7.6,"Kriti"
"Y_GE15","ES",1999,15.5,"Spain"
"Y_GE15","ES1",1999,16.5,"Noroeste (ES)"
"Y_GE15","ES11",1999,16.3,"Galicia"
"Y_GE15","ES12",1999,17.7,"Principado de Asturias"
"Y_GE15","ES13",1999,15,"Cantabria"
"Y_GE15","ES2",1999,11.6,"Noreste (ES)"
"Y_GE15","ES21",1999,14,"País Vasco"
"Y_GE15","ES22",1999,8.3,"Comunidad Foral de Navarra"
"Y_GE15","ES23",1999,6.6,"La Rioja"
"Y_GE15","ES24",1999,9.9,"Aragón"
"Y_GE15","ES3",1999,12.8,"Comunidad de Madrid"
"Y_GE15","ES30",1999,12.8,"Comunidad de Madrid"
"Y_GE15","ES4",1999,17.1,"Centro (ES)"
"Y_GE15","ES41",1999,15.2,"Castilla y León"
"Y_GE15","ES42",1999,15.1,"Castilla-la Mancha"
"Y_GE15","ES43",1999,24.9,"Extremadura"
"Y_GE15","ES5",1999,11.4,"Este (ES)"
"Y_GE15","ES51",1999,10.6,"Cataluña"
"Y_GE15","ES52",1999,13.8,"Comunidad Valenciana"
"Y_GE15","ES53",1999,7.1,"Illes Balears"
"Y_GE15","ES6",1999,24.1,"Sur (ES)"
"Y_GE15","ES61",1999,25.7,"Andalucía"
"Y_GE15","ES62",1999,14.1,"Región de Murcia"
"Y_GE15","ES63",1999,27.3,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE15","ES64",1999,21.7,"Ciudad Autónoma de Melilla (ES)"
"Y_GE15","ES7",1999,13.8,"Canarias (ES)"
"Y_GE15","ES70",1999,13.8,"Canarias (ES)"
"Y_GE15","EU15",1999,9.4,"European Union (15 countries)"
"Y_GE15","FI",1999,11.7,"Finland"
"Y_GE15","FI1",1999,11.7,"Manner-Suomi"
"Y_GE15","FI19",1999,12.8,"Länsi-Suomi"
"Y_GE15","FI2",1999,NA,"Åland"
"Y_GE15","FI20",1999,NA,"Åland"
"Y_GE15","FR",1999,12,"France"
"Y_GE15","FR1",1999,10.5,"Île de France"
"Y_GE15","FR10",1999,10.5,"Île de France"
"Y_GE15","FR2",1999,12,"Bassin Parisien"
"Y_GE15","FR21",1999,13.2,"Champagne-Ardenne"
"Y_GE15","FR22",1999,13.4,"Picardie"
"Y_GE15","FR23",1999,14.1,"Haute-Normandie"
"Y_GE15","FR24",1999,10.8,"Centre (FR)"
"Y_GE15","FR25",1999,10,"Basse-Normandie"
"Y_GE15","FR26",1999,10.4,"Bourgogne"
"Y_GE15","FR3",1999,18.1,"Nord - Pas-de-Calais"
"Y_GE15","FR30",1999,18.1,"Nord - Pas-de-Calais"
"Y_GE15","FR4",1999,9.6,"Est (FR)"
"Y_GE15","FR41",1999,11.1,"Lorraine"
"Y_GE15","FR42",1999,7.5,"Alsace"
"Y_GE15","FR43",1999,9.7,"Franche-Comté"
"Y_GE15","FR5",1999,11,"Ouest (FR)"
"Y_GE15","FR51",1999,12.2,"Pays de la Loire"
"Y_GE15","FR52",1999,9.5,"Bretagne"
"Y_GE15","FR53",1999,10.9,"Poitou-Charentes"
"Y_GE15","FR6",1999,11.3,"Sud-Ouest (FR)"
"Y_GE15","FR61",1999,11.9,"Aquitaine"
"Y_GE15","FR62",1999,11.1,"Midi-Pyrénées"
"Y_GE15","FR63",1999,9.5,"Limousin"
"Y_GE15","FR7",1999,10,"Centre-Est (FR)"
"Y_GE15","FR71",1999,9.9,"Rhône-Alpes"
"Y_GE15","FR72",1999,10.6,"Auvergne"
"Y_GE15","FR8",1999,17.4,"Méditerranée"
"Y_GE15","FR81",1999,17.4,"Languedoc-Roussillon"
"Y_GE15","FR82",1999,16.9,"Provence-Alpes-Côte d'Azur"
"Y_GE15","FR83",1999,26,"Corse"
"Y_GE15","HU",1999,6.9,"Hungary"
"Y_GE15","HU1",1999,4.9,"Közép-Magyarország"
"Y_GE15","HU10",1999,4.9,"Közép-Magyarország"
"Y_GE15","HU2",1999,6.3,"Dunántúl"
"Y_GE15","HU21",1999,6.2,"Közép-Dunántúl"
"Y_GE15","HU22",1999,4.5,"Nyugat-Dunántúl"
"Y_GE15","HU23",1999,8.4,"Dél-Dunántúl"
"Y_GE15","HU3",1999,9.1,"Alföld és Észak"
"Y_GE15","HU31",1999,11.7,"Észak-Magyarország"
"Y_GE15","HU32",1999,10,"Észak-Alföld"
"Y_GE15","HU33",1999,5.9,"Dél-Alföld"
"Y_GE15","IE",1999,5.8,"Ireland"
"Y_GE15","IE0",1999,5.8,"Éire/Ireland"
"Y_GE15","IE01",1999,6.9,"Border, Midland and Western"
"Y_GE15","IE02",1999,5.4,"Southern and Eastern"
"Y_GE15","IS",1999,2.2,"Iceland"
"Y_GE15","IS0",1999,2.2,"Ísland"
"Y_GE15","IS00",1999,2.2,"Ísland"
"Y_GE15","IT",1999,11.7,"Italy"
"Y_GE15","ITC",1999,6.2,"Nord-Ovest"
"Y_GE15","ITC1",1999,7.7,"Piemonte"
"Y_GE15","ITC2",1999,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE15","ITC3",1999,10.6,"Liguria"
"Y_GE15","ITC4",1999,4.8,"Lombardia"
"Y_GE15","ITF",1999,21.2,"Sud"
"Y_GE15","ITF1",1999,10.4,"Abruzzo"
"Y_GE15","ITF2",1999,16.3,"Molise"
"Y_GE15","ITF3",1999,23.2,"Campania"
"Y_GE15","ITF4",1999,19.5,"Puglia"
"Y_GE15","ITF5",1999,17,"Basilicata"
"Y_GE15","ITF6",1999,28.1,"Calabria"
"Y_GE15","ITG",1999,23.5,"Isole"
"Y_GE15","ITG1",1999,24.3,"Sicilia"
"Y_GE15","ITG2",1999,21.4,"Sardegna"
"Y_GE15","ITH",1999,4.8,"Nord-Est"
"Y_GE15","ITH1",1999,2.3,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE15","ITH2",1999,5.3,"Provincia Autonoma di Trento"
"Y_GE15","ITH3",1999,4.8,"Veneto"
"Y_GE15","ITH4",1999,5.5,"Friuli-Venezia Giulia"
"Y_GE15","ITI",1999,10,"Centro (IT)"
"Y_GE15","ITI1",1999,8,"Toscana"
"Y_GE15","ITI2",1999,7,"Umbria"
"Y_GE15","ITI4",1999,12.9,"Lazio"
"Y_GE15","LT",1999,13.4,"Lithuania"
"Y_GE15","LT0",1999,13.4,"Lietuva"
"Y_GE15","LT00",1999,13.4,"Lietuva"
"Y_GE15","LU",1999,2.4,"Luxembourg"
"Y_GE15","LU0",1999,2.4,"Luxembourg"
"Y_GE15","LU00",1999,2.4,"Luxembourg"
"Y_GE15","LV",1999,13.8,"Latvia"
"Y_GE15","LV0",1999,13.8,"Latvija"
"Y_GE15","LV00",1999,13.8,"Latvija"
"Y_GE15","NL",1999,3.6,"Netherlands"
"Y_GE15","NL1",1999,6.2,"Noord-Nederland"
"Y_GE15","NL11",1999,6.6,"Groningen"
"Y_GE15","NL12",1999,4.1,"Friesland (NL)"
"Y_GE15","NL13",1999,8.4,"Drenthe"
"Y_GE15","NL2",1999,3.3,"Oost-Nederland"
"Y_GE15","NL21",1999,3.1,"Overijssel"
"Y_GE15","NL22",1999,3.4,"Gelderland"
"Y_GE15","NL23",1999,4,"Flevoland"
"Y_GE15","NL3",1999,3.5,"West-Nederland"
"Y_GE15","NL31",1999,2.6,"Utrecht"
"Y_GE15","NL32",1999,3.7,"Noord-Holland"
"Y_GE15","NL33",1999,3.5,"Zuid-Holland"
"Y_GE15","NL34",1999,6,"Zeeland"
"Y_GE15","NL4",1999,2.9,"Zuid-Nederland"
"Y_GE15","NL41",1999,2.8,"Noord-Brabant"
"Y_GE15","NL42",1999,3.2,"Limburg (NL)"
"Y_GE15","NO",1999,3.2,"Norway"
"Y_GE15","NO0",1999,3.2,"Norge"
"Y_GE15","NO01",1999,2.3,"Oslo og Akershus"
"Y_GE15","NO02",1999,3.2,"Hedmark og Oppland"
"Y_GE15","NO03",1999,3.6,"Sør-Østlandet"
"Y_GE15","NO04",1999,3.4,"Agder og Rogaland"
"Y_GE15","NO05",1999,3.1,"Vestlandet"
"Y_GE15","NO06",1999,3.8,"Trøndelag"
"Y_GE15","NO07",1999,4.5,"Nord-Norge"
"Y_GE15","PL",1999,12.3,"Poland"
"Y_GE15","PL1",1999,10.9,"Region Centralny"
"Y_GE15","PL11",1999,12.2,"Lódzkie"
"Y_GE15","PL12",1999,10.2,"Mazowieckie"
"Y_GE15","PL2",1999,10.3,"Region Poludniowy"
"Y_GE15","PL21",1999,9.3,"Malopolskie"
"Y_GE15","PL22",1999,11.1,"Slaskie"
"Y_GE15","PL3",1999,12.2,"Region Wschodni"
"Y_GE15","PL31",1999,11,"Lubelskie"
"Y_GE15","PL32",1999,12.6,"Podkarpackie"
"Y_GE15","PL33",1999,13.2,"Swietokrzyskie"
"Y_GE15","PL34",1999,12.3,"Podlaskie"
"Y_GE15","PL4",1999,13.8,"Region Pólnocno-Zachodni"
"Y_GE15","PL41",1999,9.8,"Wielkopolskie"
"Y_GE15","PL42",1999,19.8,"Zachodniopomorskie"
"Y_GE15","PL43",1999,16.3,"Lubuskie"
"Y_GE15","PL5",1999,14.6,"Region Poludniowo-Zachodni"
"Y_GE15","PL51",1999,14.8,"Dolnoslaskie"
"Y_GE15","PL52",1999,14.1,"Opolskie"
"Y_GE15","PL6",1999,14,"Region Pólnocny"
"Y_GE15","PL61",1999,13.2,"Kujawsko-Pomorskie"
"Y_GE15","PL62",1999,19.5,"Warminsko-Mazurskie"
"Y_GE15","PL63",1999,11.1,"Pomorskie"
"Y_GE15","PT",1999,4.6,"Portugal"
"Y_GE15","PT1",1999,4.6,"Continente"
"Y_GE15","PT11",1999,4.6,"Norte"
"Y_GE15","PT15",1999,NA,"Algarve"
"Y_GE15","PT16",1999,2.5,"Centro (PT)"
"Y_GE15","PT17",1999,6.1,"Área Metropolitana de Lisboa"
"Y_GE15","PT18",1999,7.4,"Alentejo"
"Y_GE15","PT2",1999,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT20",1999,NA,"Região Autónoma dos Açores (PT)"
"Y_GE15","PT3",1999,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","PT30",1999,NA,"Região Autónoma da Madeira (PT)"
"Y_GE15","RO",1999,6.2,"Romania"
"Y_GE15","RO1",1999,7,"Macroregiunea unu"
"Y_GE15","RO11",1999,6.8,"Nord-Vest"
"Y_GE15","RO12",1999,7.2,"Centru"
"Y_GE15","RO2",1999,6.9,"Macroregiunea doi"
"Y_GE15","RO21",1999,6.8,"Nord-Est"
"Y_GE15","RO22",1999,7,"Sud-Est"
"Y_GE15","RO3",1999,5.8,"Macroregiunea trei"
"Y_GE15","RO31",1999,6.3,"Sud - Muntenia"
"Y_GE15","RO32",1999,4.8,"Bucuresti - Ilfov"
"Y_GE15","RO4",1999,5,"Macroregiunea patru"
"Y_GE15","RO41",1999,4,"Sud-Vest Oltenia"
"Y_GE15","RO42",1999,6.4,"Vest"
"Y_GE15","SE",1999,7.6,"Sweden"
"Y_GE15","SE1",1999,6,"Östra Sverige"
"Y_GE15","SE11",1999,3.9,"Stockholm"
"Y_GE15","SE12",1999,8.4,"Östra Mellansverige"
"Y_GE15","SE2",1999,7.7,"Södra Sverige"
"Y_GE15","SE21",1999,7.4,"Småland med öarna"
"Y_GE15","SE22",1999,8.8,"Sydsverige"
"Y_GE15","SE23",1999,7,"Västsverige"
"Y_GE15","SE3",1999,10.5,"Norra Sverige"
"Y_GE15","SE31",1999,11,"Norra Mellansverige"
"Y_GE15","SE32",1999,8.3,"Mellersta Norrland"
"Y_GE15","SE33",1999,11.5,"Övre Norrland"
"Y_GE15","SI",1999,7.3,"Slovenia"
"Y_GE15","SI0",1999,7.3,"Slovenija"
"Y_GE15","SK",1999,15.9,"Slovakia"
"Y_GE15","SK0",1999,15.9,"Slovensko"
"Y_GE15","SK01",1999,7,"Bratislavský kraj"
"Y_GE15","SK02",1999,14.1,"Západné Slovensko"
"Y_GE15","SK03",1999,18.2,"Stredné Slovensko"
"Y_GE15","SK04",1999,20.5,"Východné Slovensko"
"Y_GE15","UK",1999,6,"United Kingdom"
"Y_GE15","UKC",1999,10,"North East (UK)"
"Y_GE15","UKC1",1999,10.4,"Tees Valley and Durham"
"Y_GE15","UKC2",1999,9.8,"Northumberland and Tyne and Wear"
"Y_GE15","UKD",1999,6.2,"North West (UK)"
"Y_GE15","UKD1",1999,6.2,"Cumbria"
"Y_GE15","UKD3",1999,6.3,"Greater Manchester"
"Y_GE15","UKD4",1999,4.2,"Lancashire"
"Y_GE15","UKE",1999,6.6,"Yorkshire and The Humber"
"Y_GE15","UKE1",1999,8.6,"East Yorkshire and Northern Lincolnshire"
"Y_GE15","UKE2",1999,3.8,"North Yorkshire"
"Y_GE15","UKE3",1999,7.9,"South Yorkshire"
"Y_GE15","UKE4",1999,6,"West Yorkshire"
"Y_GE15","UKF",1999,5.2,"East Midlands (UK)"
"Y_GE15","UKF1",1999,5.7,"Derbyshire and Nottinghamshire"
"Y_GE15","UKF2",1999,4.8,"Leicestershire, Rutland and Northamptonshire"
"Y_GE15","UKF3",1999,4.7,"Lincolnshire"
"Y_GE15","UKG",1999,6.9,"West Midlands (UK)"
"Y_GE15","UKG1",1999,4.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE15","UKG2",1999,6.2,"Shropshire and Staffordshire"
"Y_GE15","UKG3",1999,8.4,"West Midlands"
"Y_GE15","UKH",1999,4.2,"East of England"
"Y_GE15","UKH1",1999,4.1,"East Anglia"
"Y_GE15","UKH2",1999,4.1,"Bedfordshire and Hertfordshire"
"Y_GE15","UKH3",1999,4.4,"Essex"
"Y_GE15","UKI",1999,7.6,"London"
"Y_GE15","UKI1",1999,9.5,"Inner London (NUTS 2010)"
"Y_GE15","UKI2",1999,6.5,"Outer London (NUTS 2010)"
"Y_GE15","UKJ",1999,3.7,"South East (UK)"
"Y_GE15","UKJ1",1999,2.6,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE15","UKJ2",1999,3.6,"Surrey, East and West Sussex"
"Y_GE15","UKJ3",1999,4.6,"Hampshire and Isle of Wight"
"Y_GE15","UKJ4",1999,4.4,"Kent"
"Y_GE15","UKK",1999,4.8,"South West (UK)"
"Y_GE15","UKK1",1999,3.3,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE15","UKK2",1999,5.1,"Dorset and Somerset"
"Y_GE15","UKK3",1999,7.7,"Cornwall and Isles of Scilly"
"Y_GE15","UKK4",1999,6.3,"Devon"
"Y_GE15","UKL",1999,7.1,"Wales"
"Y_GE15","UKL1",1999,7.5,"West Wales and The Valleys"
"Y_GE15","UKL2",1999,6.5,"East Wales"
"Y_GE15","UKM",1999,7.3,"Scotland"
"Y_GE15","UKM2",1999,6.6,"Eastern Scotland"
"Y_GE15","UKM3",1999,8.8,"South Western Scotland"
"Y_GE15","UKN",1999,7.2,"Northern Ireland (UK)"
"Y_GE15","UKN0",1999,7.2,"Northern Ireland (UK)"
"Y_GE25","AT",1999,4.5,"Austria"
"Y_GE25","AT1",1999,5.4,"Ostösterreich"
"Y_GE25","AT11",1999,4.6,"Burgenland (AT)"
"Y_GE25","AT12",1999,4.3,"Niederösterreich"
"Y_GE25","AT13",1999,6.5,"Wien"
"Y_GE25","AT2",1999,4,"Südösterreich"
"Y_GE25","AT21",1999,3.9,"Kärnten"
"Y_GE25","AT22",1999,4,"Steiermark"
"Y_GE25","AT3",1999,3.7,"Westösterreich"
"Y_GE25","AT31",1999,4.2,"Oberösterreich"
"Y_GE25","AT32",1999,3,"Salzburg"
"Y_GE25","AT33",1999,2.9,"Tirol"
"Y_GE25","AT34",1999,4,"Vorarlberg"
"Y_GE25","BE",1999,7.2,"Belgium"
"Y_GE25","BE1",1999,13.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE10",1999,13.9,"Région de Bruxelles-Capitale / Brussels Hoofdstedelijk Gewest"
"Y_GE25","BE2",1999,4.5,"Vlaams Gewest"
"Y_GE25","BE21",1999,5.4,"Prov. Antwerpen"
"Y_GE25","BE22",1999,5.6,"Prov. Limburg (BE)"
"Y_GE25","BE23",1999,5.3,"Prov. Oost-Vlaanderen"
"Y_GE25","BE24",1999,2.8,"Prov. Vlaams-Brabant"
"Y_GE25","BE25",1999,3.3,"Prov. West-Vlaanderen"
"Y_GE25","BE3",1999,10.3,"Région wallonne"
"Y_GE25","BE31",1999,6.4,"Prov. Brabant Wallon"
"Y_GE25","BE32",1999,13.9,"Prov. Hainaut"
"Y_GE25","BE33",1999,9.8,"Prov. Liège"
"Y_GE25","BE34",1999,NA,"Prov. Luxembourg (BE)"
"Y_GE25","BE35",1999,7.7,"Prov. Namur"
"Y_GE25","CH",1999,2.6,"Switzerland"
"Y_GE25","CH0",1999,2.6,"Schweiz/Suisse/Svizzera"
"Y_GE25","CZ",1999,7.2,"Czech Republic"
"Y_GE25","CZ0",1999,7.2,"Ceská republika"
"Y_GE25","CZ01",1999,3,"Praha"
"Y_GE25","CZ02",1999,7,"Strední Cechy"
"Y_GE25","CZ03",1999,5.4,"Jihozápad"
"Y_GE25","CZ04",1999,11.2,"Severozápad"
"Y_GE25","CZ05",1999,6.3,"Severovýchod"
"Y_GE25","CZ06",1999,6.8,"Jihovýchod"
"Y_GE25","CZ07",1999,8.1,"Strední Morava"
"Y_GE25","CZ08",1999,10.4,"Moravskoslezsko"
"Y_GE25","DE",1999,8.9,"Germany (until 1990 former territory of the FRG)"
"Y_GE25","DE1",1999,5.5,"Baden-Württemberg"
"Y_GE25","DE11",1999,5.4,"Stuttgart"
"Y_GE25","DE12",1999,6.3,"Karlsruhe"
"Y_GE25","DE13",1999,5.2,"Freiburg"
"Y_GE25","DE14",1999,4.7,"Tübingen"
"Y_GE25","DE2",1999,4.9,"Bayern"
"Y_GE25","DE21",1999,3.9,"Oberbayern"
"Y_GE25","DE22",1999,5.1,"Niederbayern"
"Y_GE25","DE23",1999,4.4,"Oberpfalz"
"Y_GE25","DE24",1999,6.1,"Oberfranken"
"Y_GE25","DE25",1999,6.4,"Mittelfranken"
"Y_GE25","DE26",1999,5.9,"Unterfranken"
"Y_GE25","DE27",1999,4.5,"Schwaben"
"Y_GE25","DE3",1999,15.1,"Berlin"
"Y_GE25","DE30",1999,15.1,"Berlin"
"Y_GE25","DE4",1999,16.1,"Brandenburg"
"Y_GE25","DE40",1999,16.1,"Brandenburg"
"Y_GE25","DE5",1999,11.4,"Bremen"
"Y_GE25","DE50",1999,11.4,"Bremen"
"Y_GE25","DE6",1999,8.4,"Hamburg"
"Y_GE25","DE60",1999,8.4,"Hamburg"
"Y_GE25","DE7",1999,7.1,"Hessen"
"Y_GE25","DE71",1999,6.8,"Darmstadt"
"Y_GE25","DE72",1999,7.1,"Gießen"
"Y_GE25","DE73",1999,8.4,"Kassel"
"Y_GE25","DE8",1999,19.3,"Mecklenburg-Vorpommern"
"Y_GE25","DE80",1999,19.3,"Mecklenburg-Vorpommern"
"Y_GE25","DE9",1999,7.2,"Niedersachsen"
"Y_GE25","DE91",1999,8.4,"Braunschweig"
"Y_GE25","DE92",1999,8.2,"Hannover"
"Y_GE25","DE93",1999,6.2,"Lüneburg"
"Y_GE25","DE94",1999,6.2,"Weser-Ems"
"Y_GE25","DEA",1999,7.2,"Nordrhein-Westfalen"
"Y_GE25","DEA1",1999,7.4,"Düsseldorf"
"Y_GE25","DEA2",1999,6.7,"Köln"
"Y_GE25","DEA3",1999,7,"Münster"
"Y_GE25","DEA4",1999,6.3,"Detmold"
"Y_GE25","DEA5",1999,8.1,"Arnsberg"
"Y_GE25","DEB",1999,5.9,"Rheinland-Pfalz"
"Y_GE25","DEB1",1999,5.4,"Koblenz"
"Y_GE25","DEB2",1999,5.9,"Trier"
"Y_GE25","DEB3",1999,6.3,"Rheinhessen-Pfalz"
"Y_GE25","DEC",1999,7.2,"Saarland"
"Y_GE25","DEC0",1999,7.2,"Saarland"
"Y_GE25","DED",1999,16.8,"Sachsen"
"Y_GE25","DEE",1999,21.9,"Sachsen-Anhalt"
"Y_GE25","DEE0",1999,21.9,"Sachsen-Anhalt"
"Y_GE25","DEF",1999,7.4,"Schleswig-Holstein"
"Y_GE25","DEF0",1999,7.4,"Schleswig-Holstein"
"Y_GE25","DEG",1999,15.4,"Thüringen"
"Y_GE25","DEG0",1999,15.4,"Thüringen"
"Y_GE25","DK",1999,4.3,"Denmark"
"Y_GE25","DK0",1999,4.3,"Danmark"
"Y_GE25","EE",1999,10.3,"Estonia"
"Y_GE25","EE0",1999,10.3,"Eesti"
"Y_GE25","EE00",1999,10.3,"Eesti"
"Y_GE25","EL",1999,9,"Greece"
"Y_GE25","EL1",1999,9.6,"Voreia Ellada (NUTS 2010)"
"Y_GE25","EL11",1999,10.1,"Anatoliki Makedonia, Thraki (NUTS 2010)"
"Y_GE25","EL12",1999,9.2,"Kentriki Makedonia (NUTS 2010)"
"Y_GE25","EL13",1999,10.1,"Dytiki Makedonia (NUTS 2010)"
"Y_GE25","EL14",1999,10.2,"Thessalia (NUTS 2010)"
"Y_GE25","EL2",1999,8.2,"Kentriki Ellada (NUTS 2010)"
"Y_GE25","EL21",1999,10.8,"Ipeiros (NUTS 2010)"
"Y_GE25","EL22",1999,3.9,"Ionia Nisia (NUTS 2010)"
"Y_GE25","EL23",1999,8.3,"Dytiki Ellada (NUTS 2010)"
"Y_GE25","EL24",1999,11.3,"Sterea Ellada (NUTS 2010)"
"Y_GE25","EL25",1999,5.4,"Peloponnisos (NUTS 2010)"
"Y_GE25","EL3",1999,9.8,"Attiki"
"Y_GE25","EL30",1999,9.8,"Attiki"
"Y_GE25","EL4",1999,6.2,"Nisia Aigaiou, Kriti"
"Y_GE25","EL41",1999,9.1,"Voreio Aigaio"
"Y_GE25","EL42",1999,5.9,"Notio Aigaio"
"Y_GE25","EL43",1999,5.6,"Kriti"
"Y_GE25","ES",1999,13.2,"Spain"
"Y_GE25","ES1",1999,14,"Noroeste (ES)"
"Y_GE25","ES11",1999,14.2,"Galicia"
"Y_GE25","ES12",1999,14.2,"Principado de Asturias"
"Y_GE25","ES13",1999,12.7,"Cantabria"
"Y_GE25","ES2",1999,10.1,"Noreste (ES)"
"Y_GE25","ES21",1999,12,"País Vasco"
"Y_GE25","ES22",1999,7.4,"Comunidad Foral de Navarra"
"Y_GE25","ES23",1999,5.4,"La Rioja"
"Y_GE25","ES24",1999,8.9,"Aragón"
"Y_GE25","ES3",1999,11,"Comunidad de Madrid"
"Y_GE25","ES30",1999,11,"Comunidad de Madrid"
"Y_GE25","ES4",1999,14.6,"Centro (ES)"
"Y_GE25","ES41",1999,12.8,"Castilla y León"
"Y_GE25","ES42",1999,13,"Castilla-la Mancha"
"Y_GE25","ES43",1999,21.9,"Extremadura"
"Y_GE25","ES5",1999,9.5,"Este (ES)"
"Y_GE25","ES51",1999,8.8,"Cataluña"
"Y_GE25","ES52",1999,11.5,"Comunidad Valenciana"
"Y_GE25","ES53",1999,6,"Illes Balears"
"Y_GE25","ES6",1999,21,"Sur (ES)"
"Y_GE25","ES61",1999,22.6,"Andalucía"
"Y_GE25","ES62",1999,11.5,"Región de Murcia"
"Y_GE25","ES63",1999,21.2,"Ciudad Autónoma de Ceuta (ES)"
"Y_GE25","ES64",1999,16.7,"Ciudad Autónoma de Melilla (ES)"
"Y_GE25","ES7",1999,11.1,"Canarias (ES)"
"Y_GE25","ES70",1999,11.1,"Canarias (ES)"
"Y_GE25","EU15",1999,8.2,"European Union (15 countries)"
"Y_GE25","FI",1999,8.7,"Finland"
"Y_GE25","FI1",1999,8.7,"Manner-Suomi"
"Y_GE25","FI19",1999,9.6,"Länsi-Suomi"
"Y_GE25","FI2",1999,NA,"Åland"
"Y_GE25","FI20",1999,NA,"Åland"
"Y_GE25","FR",1999,10.4,"France"
"Y_GE25","FR1",1999,9.5,"Île de France"
"Y_GE25","FR10",1999,9.5,"Île de France"
"Y_GE25","FR2",1999,10.1,"Bassin Parisien"
"Y_GE25","FR21",1999,11.2,"Champagne-Ardenne"
"Y_GE25","FR22",1999,11.1,"Picardie"
"Y_GE25","FR23",1999,11.4,"Haute-Normandie"
"Y_GE25","FR24",1999,9.6,"Centre (FR)"
"Y_GE25","FR25",1999,8.3,"Basse-Normandie"
"Y_GE25","FR26",1999,9,"Bourgogne"
"Y_GE25","FR3",1999,14.9,"Nord - Pas-de-Calais"
"Y_GE25","FR30",1999,14.9,"Nord - Pas-de-Calais"
"Y_GE25","FR4",1999,8.3,"Est (FR)"
"Y_GE25","FR41",1999,9.7,"Lorraine"
"Y_GE25","FR42",1999,6.3,"Alsace"
"Y_GE25","FR43",1999,8.4,"Franche-Comté"
"Y_GE25","FR5",1999,9.4,"Ouest (FR)"
"Y_GE25","FR51",1999,10.8,"Pays de la Loire"
"Y_GE25","FR52",1999,8.1,"Bretagne"
"Y_GE25","FR53",1999,8.8,"Poitou-Charentes"
"Y_GE25","FR6",1999,9.6,"Sud-Ouest (FR)"
"Y_GE25","FR61",1999,10.1,"Aquitaine"
"Y_GE25","FR62",1999,9.5,"Midi-Pyrénées"
"Y_GE25","FR63",1999,7.9,"Limousin"
"Y_GE25","FR7",1999,8.6,"Centre-Est (FR)"
"Y_GE25","FR71",1999,8.6,"Rhône-Alpes"
"Y_GE25","FR72",1999,8.6,"Auvergne"
"Y_GE25","FR8",1999,15.8,"Méditerranée"
"Y_GE25","FR81",1999,15.6,"Languedoc-Roussillon"
"Y_GE25","FR82",1999,15.5,"Provence-Alpes-Côte d'Azur"
"Y_GE25","FR83",1999,23.5,"Corse"
"Y_GE25","HU",1999,6,"Hungary"
"Y_GE25","HU1",1999,4.4,"Közép-Magyarország"
"Y_GE25","HU10",1999,4.4,"Közép-Magyarország"
"Y_GE25","HU2",1999,5.4,"Dunántúl"
"Y_GE25","HU21",1999,5.6,"Közép-Dunántúl"
"Y_GE25","HU22",1999,4.1,"Nyugat-Dunántúl"
"Y_GE25","HU23",1999,6.8,"Dél-Dunántúl"
"Y_GE25","HU3",1999,7.8,"Alföld és Észak"
"Y_GE25","HU31",1999,10.1,"Észak-Magyarország"
"Y_GE25","HU32",1999,8.7,"Észak-Alföld"
"Y_GE25","HU33",1999,4.8,"Dél-Alföld"
"Y_GE25","IE",1999,5.1,"Ireland"
"Y_GE25","IE0",1999,5.1,"Éire/Ireland"
"Y_GE25","IE01",1999,6.2,"Border, Midland and Western"
"Y_GE25","IE02",1999,4.8,"Southern and Eastern"
"Y_GE25","IS",1999,1.8,"Iceland"
"Y_GE25","IS0",1999,1.8,"Ísland"
"Y_GE25","IS00",1999,1.8,"Ísland"
"Y_GE25","IT",1999,9,"Italy"
"Y_GE25","ITC",1999,4.8,"Nord-Ovest"
"Y_GE25","ITC1",1999,5.9,"Piemonte"
"Y_GE25","ITC2",1999,NA,"Valle d'Aosta/Vallée d'Aoste"
"Y_GE25","ITC3",1999,8.4,"Liguria"
"Y_GE25","ITC4",1999,3.7,"Lombardia"
"Y_GE25","ITF",1999,16.1,"Sud"
"Y_GE25","ITF1",1999,8.2,"Abruzzo"
"Y_GE25","ITF2",1999,12.1,"Molise"
"Y_GE25","ITF3",1999,17.4,"Campania"
"Y_GE25","ITF4",1999,14.4,"Puglia"
"Y_GE25","ITF5",1999,12.7,"Basilicata"
"Y_GE25","ITF6",1999,23.1,"Calabria"
"Y_GE25","ITG",1999,18,"Isole"
"Y_GE25","ITG1",1999,18.5,"Sicilia"
"Y_GE25","ITG2",1999,16.7,"Sardegna"
"Y_GE25","ITH",1999,3.9,"Nord-Est"
"Y_GE25","ITH1",1999,NA,"Provincia Autonoma di Bolzano/Bozen"
"Y_GE25","ITH2",1999,4.8,"Provincia Autonoma di Trento"
"Y_GE25","ITH3",1999,3.9,"Veneto"
"Y_GE25","ITH4",1999,4.8,"Friuli-Venezia Giulia"
"Y_GE25","ITI",1999,7.8,"Centro (IT)"
"Y_GE25","ITI1",1999,6.6,"Toscana"
"Y_GE25","ITI2",1999,5.6,"Umbria"
"Y_GE25","ITI4",1999,9.8,"Lazio"
"Y_GE25","LT",1999,11.7,"Lithuania"
"Y_GE25","LT0",1999,11.7,"Lietuva"
"Y_GE25","LT00",1999,11.7,"Lietuva"
"Y_GE25","LU",1999,2,"Luxembourg"
"Y_GE25","LU0",1999,2,"Luxembourg"
"Y_GE25","LU00",1999,2,"Luxembourg"
"Y_GE25","LV",1999,12.4,"Latvia"
"Y_GE25","LV0",1999,12.4,"Latvija"
"Y_GE25","LV00",1999,12.4,"Latvija"
"Y_GE25","NL",1999,2.9,"Netherlands"
"Y_GE25","NL1",1999,4.8,"Noord-Nederland"
"Y_GE25","NL11",1999,5.1,"Groningen"
"Y_GE25","NL12",1999,2.9,"Friesland (NL)"
"Y_GE25","NL13",1999,7.1,"Drenthe"
"Y_GE25","NL2",1999,2.6,"Oost-Nederland"
"Y_GE25","NL21",1999,2.3,"Overijssel"
"Y_GE25","NL22",1999,2.6,"Gelderland"
"Y_GE25","NL23",1999,3.5,"Flevoland"
"Y_GE25","NL3",1999,2.9,"West-Nederland"
"Y_GE25","NL31",1999,2.6,"Utrecht"
"Y_GE25","NL32",1999,3,"Noord-Holland"
"Y_GE25","NL33",1999,2.6,"Zuid-Holland"
"Y_GE25","NL34",1999,5.3,"Zeeland"
"Y_GE25","NL4",1999,2.4,"Zuid-Nederland"
"Y_GE25","NL41",1999,2.2,"Noord-Brabant"
"Y_GE25","NL42",1999,2.6,"Limburg (NL)"
"Y_GE25","NO",1999,1.7,"Norway"
"Y_GE25","NO0",1999,1.7,"Norge"
"Y_GE25","NO01",1999,1.2,"Oslo og Akershus"
"Y_GE25","NO02",1999,1.4,"Hedmark og Oppland"
"Y_GE25","NO03",1999,2.2,"Sør-Østlandet"
"Y_GE25","NO04",1999,2.2,"Agder og Rogaland"
"Y_GE25","NO05",1999,1.5,"Vestlandet"
"Y_GE25","NO06",1999,2,"Trøndelag"
"Y_GE25","NO07",1999,2.1,"Nord-Norge"
"Y_GE25","PL",1999,10.1,"Poland"
"Y_GE25","PL1",1999,9.3,"Region Centralny"
"Y_GE25","PL11",1999,10.5,"Lódzkie"
"Y_GE25","PL12",1999,8.7,"Mazowieckie"
"Y_GE25","PL2",1999,8.3,"Region Poludniowy"
"Y_GE25","PL21",1999,6.6,"Malopolskie"
"Y_GE25","PL22",1999,9.6,"Slaskie"
"Y_GE25","PL3",1999,9.6,"Region Wschodni"
"Y_GE25","PL31",1999,8.5,"Lubelskie"
"Y_GE25","PL32",1999,9.3,"Podkarpackie"
"Y_GE25","PL33",1999,11,"Swietokrzyskie"
"Y_GE25","PL34",1999,10.5,"Podlaskie"
"Y_GE25","PL4",1999,11.1,"Region Pólnocno-Zachodni"
"Y_GE25","PL41",1999,7.7,"Wielkopolskie"
"Y_GE25","PL42",1999,15.3,"Zachodniopomorskie"
"Y_GE25","PL43",1999,14.7,"Lubuskie"
"Y_GE25","PL5",1999,12.2,"Region Poludniowo-Zachodni"
"Y_GE25","PL51",1999,12.3,"Dolnoslaskie"
"Y_GE25","PL52",1999,11.6,"Opolskie"
"Y_GE25","PL6",1999,12.3,"Region Pólnocny"
"Y_GE25","PL61",1999,11.1,"Kujawsko-Pomorskie"
"Y_GE25","PL62",1999,16.6,"Warminsko-Mazurskie"
"Y_GE25","PL63",1999,10.5,"Pomorskie"
"Y_GE25","PT",1999,3.9,"Portugal"
"Y_GE25","PT1",1999,3.9,"Continente"
"Y_GE25","PT11",1999,4,"Norte"
"Y_GE25","PT15",1999,NA,"Algarve"
"Y_GE25","PT16",1999,2,"Centro (PT)"
"Y_GE25","PT17",1999,5.2,"Área Metropolitana de Lisboa"
"Y_GE25","PT18",1999,6.4,"Alentejo"
"Y_GE25","PT2",1999,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT20",1999,NA,"Região Autónoma dos Açores (PT)"
"Y_GE25","PT3",1999,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","PT30",1999,NA,"Região Autónoma da Madeira (PT)"
"Y_GE25","RO",1999,4.6,"Romania"
"Y_GE25","RO1",1999,5,"Macroregiunea unu"
"Y_GE25","RO11",1999,4.9,"Nord-Vest"
"Y_GE25","RO12",1999,5.1,"Centru"
"Y_GE25","RO2",1999,5.2,"Macroregiunea doi"
"Y_GE25","RO21",1999,5.1,"Nord-Est"
"Y_GE25","RO22",1999,5.5,"Sud-Est"
"Y_GE25","RO3",1999,3.9,"Macroregiunea trei"
"Y_GE25","RO31",1999,4.3,"Sud - Muntenia"
"Y_GE25","RO32",1999,3,"Bucuresti - Ilfov"
"Y_GE25","RO4",1999,4.1,"Macroregiunea patru"
"Y_GE25","RO41",1999,3.2,"Sud-Vest Oltenia"
"Y_GE25","RO42",1999,5.3,"Vest"
"Y_GE25","SE",1999,6.7,"Sweden"
"Y_GE25","SE1",1999,5,"Östra Sverige"
"Y_GE25","SE11",1999,3.5,"Stockholm"
"Y_GE25","SE12",1999,6.9,"Östra Mellansverige"
"Y_GE25","SE2",1999,6.7,"Södra Sverige"
"Y_GE25","SE21",1999,6.7,"Småland med öarna"
"Y_GE25","SE22",1999,7.5,"Sydsverige"
"Y_GE25","SE23",1999,6.1,"Västsverige"
"Y_GE25","SE3",1999,9.7,"Norra Sverige"
"Y_GE25","SE31",1999,9.7,"Norra Mellansverige"
"Y_GE25","SE32",1999,7.7,"Mellersta Norrland"
"Y_GE25","SE33",1999,11.3,"Övre Norrland"
"Y_GE25","SI",1999,5.7,"Slovenia"
"Y_GE25","SI0",1999,5.7,"Slovenija"
"Y_GE25","SK",1999,12.8,"Slovakia"
"Y_GE25","SK0",1999,12.8,"Slovensko"
"Y_GE25","SK01",1999,5.6,"Bratislavský kraj"
"Y_GE25","SK02",1999,11.4,"Západné Slovensko"
"Y_GE25","SK03",1999,14.7,"Stredné Slovensko"
"Y_GE25","SK04",1999,16.5,"Východné Slovensko"
"Y_GE25","UK",1999,4.9,"United Kingdom"
"Y_GE25","UKC",1999,8.6,"North East (UK)"
"Y_GE25","UKC1",1999,8.8,"Tees Valley and Durham"
"Y_GE25","UKC2",1999,8.4,"Northumberland and Tyne and Wear"
"Y_GE25","UKD",1999,4.9,"North West (UK)"
"Y_GE25","UKD1",1999,5.5,"Cumbria"
"Y_GE25","UKD3",1999,4.5,"Greater Manchester"
"Y_GE25","UKD4",1999,3.4,"Lancashire"
"Y_GE25","UKE",1999,5.6,"Yorkshire and The Humber"
"Y_GE25","UKE1",1999,6.7,"East Yorkshire and Northern Lincolnshire"
"Y_GE25","UKE2",1999,NA,"North Yorkshire"
"Y_GE25","UKE3",1999,6.8,"South Yorkshire"
"Y_GE25","UKE4",1999,5.2,"West Yorkshire"
"Y_GE25","UKF",1999,3.7,"East Midlands (UK)"
"Y_GE25","UKF1",1999,4.1,"Derbyshire and Nottinghamshire"
"Y_GE25","UKF2",1999,3.4,"Leicestershire, Rutland and Northamptonshire"
"Y_GE25","UKF3",1999,NA,"Lincolnshire"
"Y_GE25","UKG",1999,5.7,"West Midlands (UK)"
"Y_GE25","UKG1",1999,3.8,"Herefordshire, Worcestershire and Warwickshire"
"Y_GE25","UKG2",1999,5,"Shropshire and Staffordshire"
"Y_GE25","UKG3",1999,7.1,"West Midlands"
"Y_GE25","UKH",1999,3.4,"East of England"
"Y_GE25","UKH1",1999,3.3,"East Anglia"
"Y_GE25","UKH2",1999,3,"Bedfordshire and Hertfordshire"
"Y_GE25","UKH3",1999,4.1,"Essex"
"Y_GE25","UKI",1999,6.5,"London"
"Y_GE25","UKI1",1999,8.3,"Inner London (NUTS 2010)"
"Y_GE25","UKI2",1999,5.5,"Outer London (NUTS 2010)"
"Y_GE25","UKJ",1999,3.1,"South East (UK)"
"Y_GE25","UKJ1",1999,2.6,"Berkshire, Buckinghamshire and Oxfordshire"
"Y_GE25","UKJ2",1999,3.2,"Surrey, East and West Sussex"
"Y_GE25","UKJ3",1999,3.5,"Hampshire and Isle of Wight"
"Y_GE25","UKJ4",1999,3.4,"Kent"
"Y_GE25","UKK",1999,3.7,"South West (UK)"
"Y_GE25","UKK1",1999,2.5,"Gloucestershire, Wiltshire and Bristol/Bath area"
"Y_GE25","UKK2",1999,4,"Dorset and Somerset"
"Y_GE25","UKK3",1999,7,"Cornwall and Isles of Scilly"
"Y_GE25","UKK4",1999,4.8,"Devon"
"Y_GE25","UKL",1999,5.3,"Wales"
"Y_GE25","UKL1",1999,5.8,"West Wales and The Valleys"
"Y_GE25","UKL2",1999,4.6,"East Wales"
"Y_GE25","UKM",1999,5.8,"Scotland"
"Y_GE25","UKM2",1999,4.8,"Eastern Scotland"
"Y_GE25","UKM3",1999,7,"South Western Scotland"
"Y_GE25","UKN",1999,6.6,"Northern Ireland (UK)"
"Y_GE25","UKN0",1999,6.6,"Northern Ireland (UK)"
